CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
7
14 Logic Display~
6 187 113 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
45199.7 5
0
14 Logic Display~
6 431 109 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
45199.7 4
0
14 Logic Display~
6 473 109 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
45199.7 3
0
9 Inverter~
13 267 203 0 2 22
0 2 3
0
0 0 608 0
6 74LS04
-21 -19 21 -11
1 S
-4 -20 3 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3670 0 0
2
45199.7 2
0
8 Hex Key~
166 147 122 0 11 12
0 2 6 7 8 0 0 0 0 0
5 53
0
0 0 4640 0
0
1 S
-4 -34 3 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
5616 0 0
2
45199.7 1
0
12 Hex Display~
7 527 124 0 18 19
10 3 2 4 5 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 M
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9323 0 0
2
45199.7 0
0
13 IAGO.Decode1b
94 302 392 0 1 7
0 0
13 IAGO.Decode1b
1 0 4736 0
0
2 U1
77 -9 91 -1
0
0
0
0
0
0
7

0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
317 0 0
2
45199.7 0
0
12
2 0 0 0 0 0 0 7 0 0 10 2
334 426
473 426
1 0 0 0 0 0 0 7 0 0 11 3
271 425
271 434
431 434
3 0 0 0 0 0 0 7 0 0 12 3
302 348
302 341
187 341
2 0 2 0 0 16 0 6 0 0 11 3
530 148
530 181
431 181
1 0 3 0 0 16 0 6 0 0 10 3
536 148
536 167
473 167
1 0 2 0 0 16 0 5 0 0 12 3
156 146
156 159
187 159
2 0 3 0 0 16 0 4 0 0 10 2
288 203
473 203
0 0 2 0 0 16 0 0 0 12 11 2
187 313
431 313
0 1 2 0 0 16 0 0 4 12 0 2
187 203
252 203
1 0 3 0 0 16 0 3 0 0 0 2
473 127
473 446
1 0 2 0 0 16 0 2 0 0 0 2
431 127
431 449
1 0 2 0 0 16 0 1 0 0 0 2
187 131
187 450
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
