CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
-1424 28 -2 779
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
-1256 124 -1143 221
9961490 0
0
6 Title:
5 Name:
0
0
0
20
13 IAGO.Decode.2
94 728 276 0 6 13
0 11 12 13 14 15 16
13 IAGO.Decode.2
3 0 4736 0
0
2 U3
74 -5 88 3
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
1 U
523 0 0
2
45190.6 18
0
14 Logic Display~
6 385 145 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
45190.6 17
0
14 Logic Display~
6 440 144 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
45190.6 16
0
14 Logic Display~
6 414 145 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
45190.6 15
0
14 Logic Display~
6 466 144 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
45190.6 14
0
8 Hex Key~
166 330 231 0 11 12
0 7 34 35 36 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I0
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
4212 0 0
2
45190.6 13
0
8 Hex Key~
166 333 317 0 11 12
0 8 31 32 33 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
4720 0 0
2
45190.6 12
0
8 Hex Key~
166 331 418 0 11 12
0 9 28 29 30 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
5551 0 0
2
45190.6 11
0
8 Hex Key~
166 332 519 0 11 12
0 10 25 26 27 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
6986 0 0
2
45190.6 10
0
8 Hex Key~
166 565 150 0 11 12
0 16 15 23 24 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 S1S0
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8745 0 0
2
45190.6 9
0
14 Logic Display~
6 604 134 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
45190.6 8
0
14 Logic Display~
6 635 133 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
45190.6 7
0
14 Logic Display~
6 916 135 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
45190.6 6
0
12 Hex Display~
7 967 143 0 16 19
10 4 20 21 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
631 0 0
2
45190.6 5
0
9 2-In AND~
219 822 376 0 3 22
0 14 7 6
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9466 0 0
2
45190.6 4
0
9 2-In AND~
219 825 426 0 3 22
0 13 8 3
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3266 0 0
2
45190.6 3
0
9 2-In AND~
219 824 480 0 3 22
0 12 9 2
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7693 0 0
2
45190.6 2
0
9 2-In AND~
219 826 531 0 3 22
0 11 10 5
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3723 0 0
2
45190.6 1
0
8 2-In OR~
219 873 449 0 3 22
0 6 5 4
0
0 0 96 0
4 4071
-15 -24 13 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3440 0 0
2
45190.6 0
0
12 IAGO.Mux.4x1
94 779 619 0 1 15
0 0
12 IAGO.Mux.4x1
1 0 4736 0
0
2 U4
71 3 85 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
6263 0 0
2
45190.6 0
0
36
5 0 0 0 0 0 0 20 0 0 33 3
812 589
812 550
466 550
6 0 0 0 0 0 0 20 0 0 34 3
786 589
786 561
440 561
4 0 0 0 0 0 0 20 0 0 35 3
759 590
759 577
414 577
3 0 0 0 0 0 0 20 0 0 36 2
728 588
385 588
2 0 0 0 0 256 0 20 0 0 27 2
701 641
604 641
1 0 0 0 0 256 0 20 0 0 26 2
701 619
635 619
7 0 0 0 0 0 0 20 0 0 32 3
779 663
779 675
916 675
3 0 2 0 0 16 0 17 0 0 0 4
845 480
855 480
855 454
866 454
3 0 3 0 0 16 0 16 0 0 0 4
846 426
854 426
854 446
867 446
1 0 4 0 0 16 0 14 0 0 32 3
976 167
976 186
916 186
3 2 5 0 0 16 0 18 19 0 0 3
847 531
860 531
860 458
3 1 6 0 0 16 0 15 19 0 0 3
843 376
860 376
860 440
3 0 4 0 0 16 0 19 0 0 32 2
906 449
916 449
2 0 7 0 0 16 0 15 0 0 33 2
798 385
466 385
2 0 8 0 0 16 0 16 0 0 34 2
801 435
440 435
2 0 9 0 0 16 0 17 0 0 35 2
800 489
414 489
2 0 10 0 0 16 0 18 0 0 36 2
802 540
385 540
1 1 11 0 0 16 0 1 18 0 0 3
678 318
678 522
802 522
2 1 12 0 0 16 0 1 17 0 0 3
700 319
700 471
800 471
3 1 13 0 0 16 0 1 16 0 0 3
728 320
728 417
801 417
4 1 14 0 0 16 0 1 15 0 0 3
762 319
762 367
798 367
0 5 15 0 0 272 0 0 1 27 0 3
604 221
679 221
679 228
0 6 16 0 0 272 0 0 1 26 0 3
635 198
760 198
760 229
2 0 15 0 0 272 0 10 0 0 27 3
568 174
568 210
604 210
1 0 16 0 0 272 0 10 0 0 26 3
574 174
574 190
635 190
1 0 16 0 0 272 0 12 0 0 0 2
635 151
635 702
1 0 15 0 0 272 0 11 0 0 0 2
604 152
604 701
1 0 10 0 0 16 0 9 0 0 36 3
341 543
341 556
385 556
1 0 9 0 0 16 0 8 0 0 35 3
340 442
340 461
414 461
1 0 8 0 0 16 0 7 0 0 34 3
342 341
342 348
440 348
1 0 7 0 0 16 0 6 0 0 33 3
339 255
339 265
466 265
1 0 4 0 0 16 0 13 0 0 0 2
916 153
916 700
1 0 7 0 0 16 0 5 0 0 0 2
466 162
466 701
1 0 8 0 0 16 0 3 0 0 0 2
440 162
440 702
1 0 9 0 0 16 0 4 0 0 0 2
414 163
414 704
1 0 10 0 0 16 0 2 0 0 0 2
385 163
385 704
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
402 78 455 102
412 86 444 102
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
538 77 591 101
548 85 580 101
4 Ctrl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
895 77 940 101
905 85 929 101
3 Out
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
