CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
11 IAGO.Add.1b
94 352 421 0 5 11
0 6 17 18 16 15
11 IAGO.Add.1b
1 0 4224 0
0
2 U1
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
4571 0 0
2
5.90093e-315 5.50185e-315
0
14 Logic Display~
6 415 147 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7796 0 0
2
5.90093e-315 5.50056e-315
0
14 Logic Display~
6 448 146 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3907 0 0
2
5.90093e-315 5.49926e-315
0
14 Logic Display~
6 478 146 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4389 0 0
2
5.90093e-315 5.49797e-315
0
14 Logic Display~
6 510 146 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7762 0 0
2
5.90093e-315 5.49667e-315
0
14 Logic Display~
6 728 145 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6723 0 0
2
5.90093e-315 5.49538e-315
0
14 Logic Display~
6 696 145 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6871 0 0
2
5.90093e-315 5.49408e-315
0
14 Logic Display~
6 666 145 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4198 0 0
2
5.90093e-315 5.49279e-315
0
14 Logic Display~
6 633 146 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
970 0 0
2
5.90093e-315 5.49149e-315
0
12 Hex Display~
7 1094 421 0 18 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 BusW
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
319 0 0
2
5.90093e-315 5.4902e-315
0
8 Hex Key~
166 373 147 0 11 12
0 8 10 13 17 0 0 0 0 0
13 68
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3663 0 0
2
5.90093e-315 5.4889e-315
0
8 Hex Key~
166 597 144 0 11 12
0 7 11 14 18 0 0 0 0 0
14 69
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3512 0 0
2
5.90093e-315 5.48761e-315
0
14 Logic Display~
6 256 404 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 Ts3
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7555 0 0
2
5.90093e-315 5.48631e-315
0
11 IAGO.Add.1b
94 541 424 0 5 11
0 5 13 14 15 12
11 IAGO.Add.1b
2 0 4224 0
0
2 U2
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
9776 0 0
2
5.90093e-315 5.46818e-315
0
11 IAGO.Add.1b
94 710 427 0 5 11
0 4 10 11 12 9
11 IAGO.Add.1b
3 0 4224 0
0
2 U3
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
6596 0 0
2
5.90093e-315 5.43451e-315
0
11 IAGO.Add.1b
94 880 430 0 5 11
0 3 8 7 9 2
11 IAGO.Add.1b
4 0 4224 0
0
2 U4
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
6750 0 0
2
5.90093e-315 5.3568e-315
0
7 Ground~
168 968 443 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9636 0 0
2
5.90093e-315 5.34643e-315
0
14 Logic Display~
6 998 407 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 W3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5369 0 0
2
5.90093e-315 5.32571e-315
0
14 Logic Display~
6 1018 406 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 W2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8555 0 0
2
5.90093e-315 5.30499e-315
0
14 Logic Display~
6 1037 405 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 W1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4690 0 0
2
5.90093e-315 5.26354e-315
0
14 Logic Display~
6 1057 403 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 W0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9145 0 0
2
5.90093e-315 0
0
11 IAGO.Add.4b
94 123 411 0 1 25
0 0
11 IAGO.Add.4b
5 0 4736 0
0
2 U5
77 1 91 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
5246 0 0
2
45187.7 0
0
68
1 0 0 0 0 0 0 22 0 0 61 2
87 456
87 545
2 0 0 0 0 0 0 22 0 0 62 2
114 456
114 526
3 0 0 0 0 0 0 22 0 0 63 2
141 455
141 510
4 0 0 0 0 0 0 22 0 0 64 2
168 455
168 491
5 0 0 0 0 0 0 22 0 0 65 2
73 378
73 253
6 0 0 0 0 0 0 22 0 0 13 2
83 378
83 234
7 0 0 0 0 0 0 22 0 0 67 2
93 378
93 218
8 0 0 0 0 0 0 22 0 0 68 2
102 378
102 199
9 0 0 0 0 0 0 22 0 0 57 2
146 378
146 343
10 0 0 0 0 0 0 22 0 0 58 2
156 377
156 324
11 0 0 0 0 0 0 22 0 0 59 2
164 377
164 308
12 0 0 0 0 0 0 22 0 0 60 2
174 378
174 289
0 0 0 0 0 0 0 0 0 66 0 2
247 234
52 234
1 0 3 0 0 4096 0 21 0 0 64 2
1057 421
1057 491
1 0 4 0 0 4096 0 20 0 0 56 2
1037 423
1037 510
1 0 5 0 0 4096 0 19 0 0 55 2
1018 424
1018 526
1 0 6 0 0 4096 0 18 0 0 61 2
998 425
998 545
3 0 7 0 0 4096 0 16 0 0 60 2
925 397
925 289
2 0 8 0 0 4096 0 16 0 0 68 2
825 397
825 199
5 1 2 0 0 8320 0 16 17 0 0 3
948 434
948 437
968 437
1 0 3 0 0 0 0 16 0 0 64 2
880 464
880 491
5 4 9 0 0 8320 0 15 16 0 0 3
778 431
778 430
803 430
2 0 10 0 0 4096 0 15 0 0 67 2
655 394
655 218
3 0 11 0 0 4096 0 15 0 0 59 2
755 394
755 308
1 0 4 0 0 0 0 15 0 0 63 2
710 461
710 510
5 4 12 0 0 8320 0 14 15 0 0 3
609 428
609 427
633 427
2 0 13 0 0 4096 0 14 0 0 66 2
486 391
486 234
3 0 14 0 0 8192 0 14 0 0 58 3
586 391
603 391
603 324
1 0 5 0 0 0 0 14 0 0 62 2
541 458
541 526
5 4 15 0 0 8320 0 1 14 0 0 3
420 425
420 424
464 424
1 4 16 0 0 8320 0 13 1 0 0 3
256 422
256 421
275 421
1 0 6 0 0 0 0 1 0 0 61 2
352 455
352 545
2 0 17 0 0 4096 0 1 0 0 65 2
297 388
297 253
3 0 18 0 0 4096 0 1 0 0 57 2
397 388
397 343
4 0 18 0 0 4096 0 12 0 0 57 2
588 168
588 343
3 0 14 0 0 4096 0 12 0 0 58 2
594 168
594 324
2 0 11 0 0 4096 0 12 0 0 59 2
600 168
600 308
1 0 7 0 0 4096 0 12 0 0 60 2
606 168
606 289
1 0 18 0 0 4096 0 9 0 0 57 2
633 164
633 343
1 0 14 0 0 4096 0 8 0 0 58 2
666 163
666 324
1 0 11 0 0 4096 0 7 0 0 59 2
696 163
696 308
1 0 7 0 0 4096 0 6 0 0 60 2
728 163
728 289
4 0 6 0 0 0 0 10 0 0 61 2
1085 445
1085 545
3 0 5 0 0 0 0 10 0 0 55 2
1091 445
1091 526
2 0 4 0 0 0 0 10 0 0 56 2
1097 445
1097 510
1 0 3 0 0 0 0 10 0 0 64 2
1103 445
1103 491
4 0 17 0 0 0 0 11 0 0 65 2
364 171
364 253
3 0 13 0 0 0 0 11 0 0 66 2
370 171
370 234
2 0 10 0 0 0 0 11 0 0 67 2
376 171
376 218
1 0 8 0 0 0 0 11 0 0 68 2
382 171
382 199
1 0 17 0 0 0 0 2 0 0 65 2
415 165
415 253
1 0 13 0 0 0 0 3 0 0 66 2
448 164
448 234
1 0 10 0 0 0 0 4 0 0 67 2
478 164
478 218
1 0 8 0 0 0 0 5 0 0 68 2
510 164
510 199
0 0 5 0 0 4096 0 0 0 62 0 2
963 526
1130 526
0 0 4 0 0 4096 0 0 0 63 0 2
959 510
1131 510
0 0 18 0 0 4224 0 0 0 0 0 2
51 343
960 343
0 0 14 0 0 4224 0 0 0 0 0 2
50 324
962 324
0 0 11 0 0 4224 0 0 0 0 0 2
50 308
958 308
0 0 7 0 0 4224 0 0 0 0 0 2
52 289
960 289
0 0 6 0 0 4224 0 0 0 0 0 2
52 545
1130 545
0 0 5 0 0 4224 0 0 0 0 0 2
53 526
967 526
0 0 4 0 0 4224 0 0 0 0 0 2
52 510
963 510
0 0 3 0 0 4224 0 0 0 0 0 2
50 491
1132 491
0 0 17 0 0 4224 0 0 0 0 0 2
48 253
953 253
0 0 13 0 0 4224 0 0 0 0 0 2
243 234
955 234
0 0 10 0 0 4224 0 0 0 0 0 2
51 218
951 218
0 0 8 0 0 4224 0 0 0 0 0 2
55 199
953 199
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1021 343 1082 367
1031 351 1071 367
5 OUT's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
506 74 559 98
516 82 548 98
4 IN's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
