CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
14
9 2-In AND~
219 334 409 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3835 0 0
2
45187.8 0
0
9 2-In AND~
219 334 359 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3670 0 0
2
45187.8 0
0
9 2-In AND~
219 334 305 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5616 0 0
2
45187.8 0
0
9 2-In AND~
219 336 256 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
45187.8 0
0
9 Inverter~
13 279 186 0 1 22
0 0
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
317 0 0
2
45187.8 0
0
9 Inverter~
13 252 186 0 1 22
0 0
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
45187.8 0
0
14 Logic Display~
6 496 112 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
45187.8 0
0
14 Logic Display~
6 522 111 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45187.8 0
0
14 Logic Display~
6 550 111 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
45187.8 0
0
14 Logic Display~
6 577 112 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
45187.8 2
0
12 Hex Display~
7 628 119 0 16 19
10 0 0 0 0 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 N3N0
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9172 0 0
2
45187.8 0
0
8 Hex Key~
166 135 110 0 11 12
0 0 0 0 0 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 S1S0
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7100 0 0
2
45187.8 0
0
14 Logic Display~
6 212 108 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
45187.8 0
0
14 Logic Display~
6 183 109 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7678 0 0
2
45187.8 0
0
29
0 0 0 0 0 256 0 0 0 0 19 5
156 158
156 637
604 637
604 143
153 143
3 0 0 0 0 0 0 1 0 0 27 2
355 409
496 409
3 0 0 0 0 0 0 2 0 0 26 2
355 359
522 359
3 0 0 0 0 0 0 3 0 0 25 2
355 305
550 305
3 0 0 0 0 0 0 4 0 0 24 2
357 256
577 256
2 0 0 0 0 256 0 2 0 0 10 2
310 368
282 368
2 0 0 0 0 256 0 4 0 0 10 2
312 265
282 265
1 0 0 0 0 256 0 4 0 0 11 2
312 247
255 247
1 0 0 0 0 0 0 3 0 0 11 2
310 296
255 296
2 0 0 0 0 256 0 5 0 0 0 2
282 204
282 610
2 0 0 0 0 256 0 6 0 0 0 2
255 204
255 608
2 0 0 0 0 0 0 3 0 0 28 2
310 314
212 314
1 0 0 0 0 0 0 2 0 0 29 2
310 350
183 350
2 0 0 0 0 0 0 1 0 0 28 2
310 418
212 418
1 0 0 0 0 0 0 1 0 0 29 2
310 400
183 400
0 1 0 0 0 0 0 0 5 28 0 3
212 130
282 130
282 168
0 1 0 0 0 0 0 0 6 29 0 3
183 137
255 137
255 168
2 0 0 0 0 0 0 12 0 0 29 3
138 134
138 150
183 150
1 0 0 0 0 0 0 12 0 0 28 3
144 134
144 143
212 143
1 0 0 0 0 0 0 11 0 0 24 3
637 143
637 181
577 181
2 0 0 0 0 0 0 11 0 0 25 3
631 143
631 171
550 171
3 0 0 0 0 0 0 11 0 0 26 3
625 143
625 163
522 163
4 0 0 0 0 0 0 11 0 0 27 3
619 143
619 157
496 157
1 0 0 0 0 0 0 10 0 0 0 2
577 130
577 611
1 0 0 0 0 0 0 9 0 0 0 2
550 129
550 612
1 0 0 0 0 0 0 8 0 0 0 2
522 129
522 614
1 0 0 0 0 0 0 7 0 0 0 2
496 130
496 614
1 0 0 0 0 0 0 13 0 0 0 2
212 126
212 613
1 0 0 0 0 0 0 14 0 0 0 2
183 127
183 614
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
346 117 439 141
356 125 428 141
9 Decode.2b
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
