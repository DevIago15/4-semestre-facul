CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
11 IAGO.Sub.1b
94 908 446 0 5 11
0 14 7 3 11 2
11 IAGO.Sub.1b
1 0 4224 0
0
2 U4
74 -44 88 -36
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
3504 0 0
2
5.90093e-315 0
0
11 IAGO.Sub.1b
94 744 443 0 5 11
0 15 8 4 12 11
11 IAGO.Sub.1b
2 0 4224 0
0
2 U3
74 -44 88 -36
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
331 0 0
2
5.90093e-315 0
0
11 IAGO.Sub.1b
94 588 440 0 5 11
0 16 9 5 13 12
11 IAGO.Sub.1b
3 0 4224 0
0
2 U2
74 -44 88 -36
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
3471 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 487 160 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5437 0 0
2
5.90093e-315 5.50056e-315
0
14 Logic Display~
6 520 159 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3177 0 0
2
5.90093e-315 5.49926e-315
0
14 Logic Display~
6 550 159 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8977 0 0
2
5.90093e-315 5.49797e-315
0
14 Logic Display~
6 582 159 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5822 0 0
2
5.90093e-315 5.49667e-315
0
14 Logic Display~
6 800 158 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5959 0 0
2
5.90093e-315 5.49538e-315
0
14 Logic Display~
6 768 158 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6537 0 0
2
5.90093e-315 5.49408e-315
0
14 Logic Display~
6 738 158 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4325 0 0
2
5.90093e-315 5.49279e-315
0
14 Logic Display~
6 705 159 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
565 0 0
2
5.90093e-315 5.49149e-315
0
12 Hex Display~
7 1166 434 0 16 19
10 14 15 16 17 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 BusZ
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3181 0 0
2
5.90093e-315 5.4902e-315
0
8 Hex Key~
166 445 160 0 11 12
0 7 8 9 10 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3758 0 0
2
5.90093e-315 5.4889e-315
0
8 Hex Key~
166 669 157 0 11 12
0 3 4 5 6 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5736 0 0
2
5.90093e-315 5.48761e-315
0
14 Logic Display~
6 328 417 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 Ts3
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6775 0 0
2
5.90093e-315 5.48631e-315
0
7 Ground~
168 1040 456 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3110 0 0
2
5.90093e-315 5.34643e-315
0
14 Logic Display~
6 1070 420 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Z3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3322 0 0
2
5.90093e-315 5.32571e-315
0
14 Logic Display~
6 1090 419 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Z2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5890 0 0
2
5.90093e-315 5.30499e-315
0
14 Logic Display~
6 1109 418 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Z1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
550 0 0
2
5.90093e-315 5.26354e-315
0
14 Logic Display~
6 1129 416 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Z0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3729 0 0
2
5.90093e-315 0
0
11 IAGO.Sub.1b
94 428 437 0 5 11
0 17 10 6 18 13
11 IAGO.Sub.1b
4 0 4224 0
0
2 U1
74 -44 88 -36
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
556 0 0
2
5.90093e-315 0
0
11 IAGO.Sub.4b
94 168 423 0 1 25
0 0
11 IAGO.Sub.4b
5 0 4736 0
0
2 U5
80 2 94 10
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3829 0 0
2
45187.7 0
0
67
5 0 0 0 0 0 0 22 0 0 64 2
115 389
115 266
6 0 0 0 0 0 0 22 0 0 65 2
128 390
128 247
7 0 0 0 0 0 0 22 0 0 66 2
141 389
141 231
8 0 0 0 0 0 0 22 0 0 67 2
150 389
150 212
9 0 0 0 0 0 0 22 0 0 56 2
195 389
195 356
10 0 0 0 0 0 0 22 0 0 57 2
204 389
204 337
11 0 0 0 0 0 0 22 0 0 58 2
213 388
213 321
12 0 0 0 0 0 0 22 0 0 59 2
223 389
223 302
1 0 0 0 0 0 0 22 0 0 60 2
132 469
132 558
2 0 0 0 0 0 0 22 0 0 61 2
159 467
159 539
3 0 0 0 0 0 0 22 0 0 62 2
186 469
186 523
4 0 0 0 0 0 0 22 0 0 63 2
214 468
214 504
3 0 3 0 0 4096 0 1 0 0 59 2
944 408
944 302
3 0 4 0 0 4096 0 2 0 0 58 2
780 405
780 321
3 0 5 0 0 4096 0 3 0 0 57 2
624 402
624 337
3 0 6 0 0 4096 0 21 0 0 56 2
464 399
464 356
2 0 7 0 0 4096 0 1 0 0 67 2
863 408
863 212
2 0 8 0 0 4096 0 2 0 0 66 2
699 405
699 231
2 0 9 0 0 4096 0 3 0 0 65 2
543 402
543 247
2 0 10 0 0 4096 0 21 0 0 64 2
383 399
383 266
5 4 11 0 0 4224 0 2 1 0 0 2
815 443
829 443
5 4 12 0 0 4224 0 3 2 0 0 2
659 440
665 440
5 4 13 0 0 4224 0 21 3 0 0 2
499 437
509 437
1 0 14 0 0 4096 0 1 0 0 63 2
908 484
908 504
1 0 15 0 0 4096 0 2 0 0 62 2
744 481
744 523
1 0 16 0 0 4096 0 3 0 0 61 2
588 478
588 539
1 0 17 0 0 4096 0 21 0 0 60 2
428 475
428 558
1 0 14 0 0 4096 0 20 0 0 63 2
1129 434
1129 504
1 0 15 0 0 4096 0 19 0 0 55 2
1109 436
1109 523
1 0 16 0 0 4096 0 18 0 0 54 2
1090 437
1090 539
1 0 17 0 0 4096 0 17 0 0 60 2
1070 438
1070 558
5 1 2 0 0 8320 0 1 16 0 0 5
979 446
979 447
1020 447
1020 450
1040 450
1 4 18 0 0 8320 0 15 21 0 0 3
328 435
328 434
349 434
4 0 6 0 0 4096 0 14 0 0 56 2
660 181
660 356
3 0 5 0 0 4096 0 14 0 0 57 2
666 181
666 337
2 0 4 0 0 4096 0 14 0 0 58 2
672 181
672 321
1 0 3 0 0 4096 0 14 0 0 59 2
678 181
678 302
1 0 6 0 0 4096 0 11 0 0 56 2
705 177
705 356
1 0 5 0 0 4096 0 10 0 0 57 2
738 176
738 337
1 0 4 0 0 4096 0 9 0 0 58 2
768 176
768 321
1 0 3 0 0 4096 0 8 0 0 59 2
800 176
800 302
4 0 17 0 0 0 0 12 0 0 60 2
1157 458
1157 558
3 0 16 0 0 0 0 12 0 0 54 2
1163 458
1163 539
2 0 15 0 0 0 0 12 0 0 55 2
1169 458
1169 523
1 0 14 0 0 0 0 12 0 0 63 2
1175 458
1175 504
4 0 10 0 0 0 0 13 0 0 64 2
436 184
436 266
3 0 9 0 0 0 0 13 0 0 65 2
442 184
442 247
2 0 8 0 0 0 0 13 0 0 66 2
448 184
448 231
1 0 7 0 0 0 0 13 0 0 67 2
454 184
454 212
1 0 10 0 0 0 0 4 0 0 64 2
487 178
487 266
1 0 9 0 0 0 0 5 0 0 65 2
520 177
520 247
1 0 8 0 0 0 0 6 0 0 66 2
550 177
550 231
1 0 7 0 0 0 0 7 0 0 67 2
582 177
582 212
0 0 16 0 0 4096 0 0 0 61 0 2
1035 539
1202 539
0 0 15 0 0 4096 0 0 0 62 0 2
1031 523
1203 523
0 0 6 0 0 4224 0 0 0 0 0 2
77 356
1032 356
0 0 5 0 0 4224 0 0 0 0 0 2
78 337
1034 337
0 0 4 0 0 4224 0 0 0 0 0 2
81 321
1030 321
0 0 3 0 0 4224 0 0 0 0 0 2
78 302
1032 302
0 0 17 0 0 4224 0 0 0 0 0 2
78 558
1202 558
0 0 16 0 0 4224 0 0 0 0 0 2
78 539
1039 539
0 0 15 0 0 4224 0 0 0 0 0 2
77 523
1035 523
0 0 14 0 0 4224 0 0 0 0 0 2
79 504
1204 504
0 0 10 0 0 4224 0 0 0 0 0 2
76 266
1025 266
0 0 9 0 0 4224 0 0 0 0 0 2
73 247
1027 247
0 0 8 0 0 4224 0 0 0 0 0 2
75 231
1023 231
0 0 7 0 0 4224 0 0 0 0 0 2
77 212
1025 212
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
578 87 631 111
588 95 620 111
4 IN's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1093 356 1154 380
1103 364 1143 380
5 OUT's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
