CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
14
8 Hex Key~
166 109 139 0 11 12
0 8 7 6 5 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
34 0 0
2
5.90093e-315 0
0
12 Hex Display~
7 622 310 0 18 19
10 12 11 10 9 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusX
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6357 0 0
2
45185.9 0
0
9 Inverter~
13 355 316 0 2 22
0 8 12
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
319 0 0
2
45185.9 1
0
9 Inverter~
13 324 316 0 2 22
0 7 11
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3976 0 0
2
45185.9 2
0
9 Inverter~
13 293 316 0 2 22
0 6 10
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7634 0 0
2
45185.9 3
0
9 Inverter~
13 263 317 0 2 22
0 5 9
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
523 0 0
2
45185.9 4
0
14 Logic Display~
6 478 297 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
45185.9 5
0
14 Logic Display~
6 512 296 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
45185.9 6
0
14 Logic Display~
6 544 295 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
45185.9 7
0
14 Logic Display~
6 575 296 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
45185.9 8
0
14 Logic Display~
6 253 128 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
45185.9 9
0
14 Logic Display~
6 222 127 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
45185.9 10
0
14 Logic Display~
6 190 128 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
45185.9 11
0
14 Logic Display~
6 156 129 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
45185.9 12
0
35
0 0 2 0 0 8592 0 0 0 0 0 5
257 169
399 169
399 464
251 464
251 370
0 0 3 0 0 8576 0 0 0 0 0 5
640 350
707 350
707 445
642 445
642 351
0 0 4 0 0 8576 0 0 0 0 0 5
26 177
93 177
93 272
28 272
28 178
4 0 5 0 0 4096 0 1 0 0 32 2
100 163
100 267
3 0 6 0 0 4096 0 1 0 0 33 2
106 163
106 238
2 0 7 0 0 4096 0 1 0 0 34 2
112 163
112 214
1 0 8 0 0 4096 0 1 0 0 35 2
118 163
118 193
4 0 9 0 0 4096 0 2 0 0 24 2
613 334
613 437
3 0 10 0 0 4096 0 2 0 0 25 2
619 334
619 410
2 0 11 0 0 4096 0 2 0 0 26 2
625 334
625 382
1 0 12 0 0 4096 0 2 0 0 27 2
631 334
631 358
2 0 9 0 0 0 0 6 0 0 24 2
266 335
266 437
0 1 5 0 0 0 0 0 6 32 0 3
265 267
266 267
266 299
2 0 10 0 0 0 0 5 0 0 25 2
296 334
296 410
0 1 6 0 0 0 0 0 5 33 0 3
298 238
296 238
296 298
2 0 11 0 0 0 0 4 0 0 26 2
327 334
327 382
0 1 7 0 0 8192 0 0 4 34 0 3
325 214
327 214
327 298
2 0 12 0 0 0 0 3 0 0 27 2
358 334
358 358
0 1 8 0 0 8192 0 0 3 35 0 3
356 193
358 193
358 298
1 0 9 0 0 4096 0 7 0 0 24 2
478 315
478 437
1 0 10 0 0 4096 0 8 0 0 25 2
512 314
512 410
1 0 11 0 0 4096 0 9 0 0 26 2
544 313
544 382
1 0 12 0 0 4096 0 10 0 0 27 2
575 314
575 358
0 0 9 0 0 4224 0 0 0 0 0 2
85 437
669 437
0 0 10 0 0 4224 0 0 0 0 0 2
83 410
669 410
0 0 11 0 0 4224 0 0 0 0 0 2
81 382
669 382
0 0 12 0 0 4224 0 0 0 0 0 2
78 358
669 358
1 0 5 0 0 4096 0 14 0 0 32 2
156 147
156 267
1 0 6 0 0 4096 0 13 0 0 33 2
190 146
190 238
1 0 7 0 0 0 0 12 0 0 34 2
222 145
222 214
1 0 8 0 0 0 0 11 0 0 35 2
253 146
253 193
0 0 5 0 0 4224 0 0 0 0 0 2
74 267
427 267
0 0 6 0 0 4224 0 0 0 0 0 2
71 238
427 238
0 0 7 0 0 4224 0 0 0 0 0 2
68 214
426 214
0 0 8 0 0 4224 0 0 0 0 0 2
66 193
428 193
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
292 139 393 163
302 147 382 163
10 Buffer.4b.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
649 321 702 345
659 329 691 345
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
33 149 86 173
43 157 75 173
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
537 231 598 255
547 239 587 255
5 OUT'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
158 64 211 88
168 72 200 88
4 IN'S
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
