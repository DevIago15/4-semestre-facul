CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
42991634 0
0
6 Title:
5 Name:
0
0
0
12
12 Hex Display~
7 748 150 0 18 19
10 3 2 10 11 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
3 TsZ
-11 -38 10 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8546 0 0
2
45187.7 11
0
8 Hex Key~
166 298 141 0 11 12
0 6 5 4 12 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 ABTe
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8607 0 0
2
45187.7 10
0
8 2-In OR~
219 604 319 0 3 22
0 8 7 2
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 O1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5781 0 0
2
45187.7 9
0
9 2-In AND~
219 519 280 0 3 22
0 9 6 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 AN1B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6991 0 0
2
45187.7 8
0
9 2-In AND~
219 432 323 0 3 22
0 4 5 7
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 AN1A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9631 0 0
2
45187.7 7
0
9 2-In XOR~
219 518 199 0 3 22
0 6 9 3
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 XO1B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8381 0 0
2
45187.7 6
0
14 Logic Display~
6 686 121 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Z
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6697 0 0
2
45187.7 5
0
14 Logic Display~
6 665 122 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3463 0 0
2
45187.7 4
0
9 2-In XOR~
219 427 242 0 3 22
0 4 5 9
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 XO1A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9605 0 0
2
45187.7 3
0
14 Logic Display~
6 395 122 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
936 0 0
2
45187.7 2
0
14 Logic Display~
6 375 121 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9813 0 0
2
45187.7 1
0
14 Logic Display~
6 355 121 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5286 0 0
2
45187.7 0
0
24
2 0 2 0 0 8208 0 1 0 0 21 3
751 174
751 187
665 187
1 0 3 0 0 8208 0 1 0 0 20 3
757 174
757 179
686 179
3 0 4 0 0 8208 0 2 0 0 24 3
295 165
295 187
355 187
2 0 5 0 0 8208 0 2 0 0 23 3
301 165
301 177
375 177
1 0 6 0 0 4112 0 2 0 0 22 2
307 165
395 165
0 0 4 0 0 4496 0 0 0 0 0 6
339 143
699 143
699 363
341 363
341 143
343 143
3 2 7 0 0 4240 0 5 3 0 0 4
453 323
555 323
555 328
591 328
3 0 2 0 0 16 0 3 0 0 21 2
637 319
665 319
3 1 8 0 0 4240 0 4 3 0 0 4
540 280
571 280
571 310
591 310
2 0 6 0 0 4112 0 4 0 0 22 2
495 289
395 289
1 0 9 0 0 4112 0 4 0 0 12 2
495 271
473 271
0 0 9 0 0 4368 0 0 0 17 0 2
473 242
473 275
2 0 5 0 0 16 0 5 0 0 23 2
408 332
375 332
1 0 4 0 0 16 0 5 0 0 24 2
408 314
355 314
3 0 3 0 0 4112 0 6 0 0 20 2
551 199
686 199
1 0 6 0 0 4112 0 6 0 0 22 2
502 190
395 190
3 2 9 0 0 8336 0 9 6 0 0 4
460 242
475 242
475 208
502 208
2 0 5 0 0 16 0 9 0 0 23 2
411 251
375 251
1 0 4 0 0 16 0 9 0 0 24 2
411 233
355 233
1 0 3 0 0 4240 0 7 0 0 0 2
686 139
686 364
1 0 2 0 0 4240 0 8 0 0 0 2
665 140
665 364
1 0 6 0 0 4240 0 10 0 0 0 2
395 140
395 364
1 0 5 0 0 4240 0 11 0 0 0 2
375 139
375 364
1 0 4 0 0 16 0 12 0 0 6 2
355 139
355 363
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
593 141 630 165
603 149 619 165
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
521 140 558 164
531 148 547 164
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
424 138 461 162
434 146 450 162
2 L1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
