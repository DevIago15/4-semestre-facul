CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
9961490 0
0
6 Title:
5 Name:
0
0
0
13
14 Logic Display~
6 411 171 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7130 0 0
2
45187.7 11
0
14 Logic Display~
6 431 171 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4115 0 0
2
45187.7 10
0
14 Logic Display~
6 451 172 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3197 0 0
2
45187.7 9
0
9 2-In XOR~
219 483 292 0 3 22
0 4 5 9
0
0 0 96 0
6 74LS86
-21 -24 21 -16
4 XO1B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
813 0 0
2
45187.7 8
0
14 Logic Display~
6 721 172 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3396 0 0
2
45187.7 7
0
14 Logic Display~
6 742 171 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Z
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6348 0 0
2
45187.7 6
0
9 2-In XOR~
219 574 249 0 3 22
0 6 9 3
0
0 0 96 0
6 74LS86
-21 -24 21 -16
4 XO1A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
583 0 0
2
45187.7 5
0
9 2-In AND~
219 488 373 0 3 22
0 4 5 7
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 AN1B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
922 0 0
2
45187.7 4
0
9 2-In AND~
219 575 330 0 3 22
0 9 6 8
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 AN1A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4442 0 0
2
45187.7 3
0
8 2-In OR~
219 660 369 0 3 22
0 8 7 2
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 O1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5893 0 0
2
45187.7 2
0
8 Hex Key~
166 354 191 0 11 12
0 6 5 4 12 0 0 0 0 0
6 54
0
0 0 4640 0
0
4 ABTe
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3814 0 0
2
45187.7 1
0
12 Hex Display~
7 804 200 0 18 19
10 3 2 10 11 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
3 TsZ
-11 -38 10 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3637 0 0
2
45187.7 0
0
11 IAGO.Sub.1b
94 585 522 0 1 11
0 0
11 IAGO.Sub.1b
1 0 4224 0
0
2 U1
74 -44 88 -36
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
6890 0 0
2
45187.7 0
0
32
4 0 0 0 0 0 0 13 0 0 29 4
506 519
495 519
495 626
721 626
1 0 0 0 0 0 0 13 0 0 28 3
585 560
585 582
742 582
0 5 0 0 0 0 0 0 13 8 0 4
451 467
662 467
662 522
656 522
0 3 0 0 0 0 0 0 13 7 0 3
431 471
621 471
621 484
2 0 0 0 0 0 0 13 0 0 6 3
540 484
540 475
411 475
0 0 0 0 0 0 0 0 0 32 0 2
411 407
411 632
0 0 0 0 0 0 0 0 0 31 0 2
431 409
431 632
0 0 0 0 0 0 0 0 0 30 0 2
451 409
451 633
2 0 2 0 0 16 0 12 0 0 29 3
807 224
807 237
721 237
1 0 3 0 0 16 0 12 0 0 28 3
813 224
813 229
742 229
3 0 4 0 0 16 0 11 0 0 32 3
351 215
351 237
411 237
2 0 5 0 0 16 0 11 0 0 31 3
357 215
357 227
431 227
1 0 6 0 0 16 0 11 0 0 30 2
363 215
451 215
0 0 4 0 0 272 0 0 0 0 0 6
395 193
755 193
755 413
397 413
397 193
399 193
3 2 7 0 0 16 0 8 10 0 0 4
509 373
611 373
611 378
647 378
3 0 2 0 0 16 0 10 0 0 29 2
693 369
721 369
3 1 8 0 0 16 0 9 10 0 0 4
596 330
627 330
627 360
647 360
2 0 6 0 0 16 0 9 0 0 30 2
551 339
451 339
1 0 9 0 0 16 0 9 0 0 20 2
551 321
529 321
0 0 9 0 0 272 0 0 0 25 0 2
529 292
529 325
2 0 5 0 0 16 0 8 0 0 31 2
464 382
431 382
1 0 4 0 0 16 0 8 0 0 32 2
464 364
411 364
3 0 3 0 0 16 0 7 0 0 28 2
607 249
742 249
1 0 6 0 0 16 0 7 0 0 30 2
558 240
451 240
3 2 9 0 0 16 0 4 7 0 0 4
516 292
531 292
531 258
558 258
2 0 5 0 0 16 0 4 0 0 31 2
467 301
431 301
1 0 4 0 0 16 0 4 0 0 32 2
467 283
411 283
1 0 3 0 0 16 0 6 0 0 0 2
742 189
742 635
1 0 2 0 0 16 0 5 0 0 0 2
721 190
721 636
1 0 6 0 0 16 0 3 0 0 0 2
451 190
451 414
1 0 5 0 0 16 0 2 0 0 0 2
431 189
431 414
1 0 4 0 0 16 0 1 0 0 14 2
411 189
411 413
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
649 191 686 215
659 199 675 215
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
577 190 614 214
587 198 603 214
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
480 188 517 212
490 196 506 212
2 L1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
