CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
12
12 Hex Display~
7 587 165 0 18 19
10 3 2 11 12 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
7 DECIMAL
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3536 0 0
2
45168.9 0
0
8 Hex Key~
166 137 156 0 11 12
0 6 5 4 13 0 0 0 0 0
7 55
0
0 0 4656 0
0
6 SOURCE
-21 -34 21 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
4597 0 0
2
45168.9 0
0
8 2-In OR~
219 443 334 0 3 22
0 9 8 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
45168.9 0
0
9 2-In AND~
219 358 295 0 3 22
0 10 6 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3670 0 0
2
45168.9 0
0
9 2-In AND~
219 271 338 0 3 22
0 4 5 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5616 0 0
2
45168.9 0
0
9 2-In XOR~
219 357 214 0 3 22
0 6 10 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOB
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
45168.9 0
0
14 Logic Display~
6 525 136 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 W
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
45168.9 1
0
14 Logic Display~
6 504 137 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45168.9 0
0
9 2-In XOR~
219 266 257 0 3 22
0 4 5 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4299 0 0
2
45168.9 0
0
14 Logic Display~
6 234 137 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
45168.9 0
0
14 Logic Display~
6 214 136 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
45168.9 0
0
14 Logic Display~
6 194 136 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
45168.9 0
0
24
2 0 2 0 0 8192 0 1 0 0 21 3
590 189
590 202
504 202
1 0 3 0 0 8192 0 1 0 0 20 3
596 189
596 194
525 194
3 0 4 0 0 8192 0 2 0 0 24 3
134 180
134 202
194 202
2 0 5 0 0 8192 0 2 0 0 23 3
140 180
140 192
214 192
1 0 6 0 0 4096 0 2 0 0 22 2
146 180
234 180
0 0 7 0 0 4480 0 0 0 0 0 6
178 158
538 158
538 378
180 378
180 158
182 158
3 2 8 0 0 4224 0 5 3 0 0 4
292 338
394 338
394 343
430 343
3 0 2 0 0 0 0 3 0 0 21 2
476 334
504 334
3 1 9 0 0 4224 0 4 3 0 0 4
379 295
410 295
410 325
430 325
2 0 6 0 0 4096 0 4 0 0 22 2
334 304
234 304
1 0 10 0 0 4096 0 4 0 0 12 2
334 286
312 286
0 0 10 0 0 4352 0 0 0 17 0 2
312 257
312 290
2 0 5 0 0 0 0 5 0 0 23 2
247 347
214 347
1 0 4 0 0 0 0 5 0 0 24 2
247 329
194 329
3 0 3 0 0 4096 0 6 0 0 20 2
390 214
525 214
1 0 6 0 0 4096 0 6 0 0 22 2
341 205
234 205
3 2 10 0 0 8320 0 9 6 0 0 4
299 257
314 257
314 223
341 223
2 0 5 0 0 0 0 9 0 0 23 2
250 266
214 266
1 0 4 0 0 0 0 9 0 0 24 2
250 248
194 248
1 0 3 0 0 4224 0 7 0 0 0 2
525 154
525 379
1 0 2 0 0 4224 0 8 0 0 0 2
504 155
504 379
1 0 6 0 0 4224 0 10 0 0 0 2
234 155
234 379
1 0 5 0 0 4224 0 11 0 0 0 2
214 154
214 379
1 0 4 0 0 4224 0 12 0 0 0 2
194 154
194 379
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
413 321 442 345
423 329 431 345
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
408 302 433 326
416 310 424 326
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
368 274 393 298
376 282 384 298
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
432 156 469 180
442 164 458 180
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
312 261 349 285
322 269 338 285
2 Te
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
311 178 348 202
321 186 337 202
2 Te
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
280 311 309 335
290 319 298 335
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
228 325 257 349
238 333 246 349
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 302 258 326
239 310 247 326
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
235 242 264 266
245 250 253 266
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
232 223 261 247
242 231 250 247
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
472 188 501 212
482 196 490 212
1 W
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
311 200 340 224
321 208 329 224
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
375 187 404 211
385 195 393 211
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
285 232 314 256
295 240 303 256
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
360 155 397 179
370 163 386 179
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 153 300 177
273 161 289 177
2 L1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
