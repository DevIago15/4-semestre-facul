CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
9961490 0
0
6 Title:
5 Name:
0
0
0
20
9 2-In AND~
219 972 469 0 3 22
0 13 9 5
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 A1D
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3138 0 0
2
5.90093e-315 5.43451e-315
0
9 2-In AND~
219 920 468 0 3 22
0 12 8 4
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 A1C
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5409 0 0
2
5.90093e-315 5.43192e-315
0
9 2-In AND~
219 872 468 0 3 22
0 11 7 3
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 A1B
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
983 0 0
2
5.90093e-315 5.42933e-315
0
9 2-In AND~
219 822 470 0 3 22
0 10 6 2
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 A1A
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6652 0 0
2
5.90093e-315 5.42414e-315
0
14 Logic Display~
6 718 210 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4281 0 0
2
5.90093e-315 5.41896e-315
0
14 Logic Display~
6 684 209 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6847 0 0
2
5.90093e-315 5.41378e-315
0
14 Logic Display~
6 646 210 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6543 0 0
2
5.90093e-315 5.4086e-315
0
14 Logic Display~
6 608 210 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90093e-315 5.40342e-315
0
8 Hex Key~
166 557 213 0 11 12
0 13 12 11 10 0 0 0 0 0
14 69
0
0 0 4656 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3828 0 0
2
5.90093e-315 5.39824e-315
0
14 Logic Display~
6 1128 460 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
955 0 0
2
5.90093e-315 5.39306e-315
0
14 Logic Display~
6 1097 459 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7782 0 0
2
5.90093e-315 5.38788e-315
0
14 Logic Display~
6 1065 460 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
824 0 0
2
5.90093e-315 5.37752e-315
0
14 Logic Display~
6 1031 461 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6983 0 0
2
5.90093e-315 5.36716e-315
0
12 Hex Display~
7 1175 474 0 18 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusY
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3185 0 0
2
5.90093e-315 5.3568e-315
0
8 Hex Key~
166 350 220 0 11 12
0 9 8 7 6 0 0 0 0 0
10 65
0
0 0 4656 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4213 0 0
2
5.90093e-315 5.34643e-315
0
14 Logic Display~
6 494 209 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9765 0 0
2
5.90093e-315 5.32571e-315
0
14 Logic Display~
6 463 208 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8986 0 0
2
5.90093e-315 5.30499e-315
0
14 Logic Display~
6 431 209 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3273 0 0
2
5.90093e-315 5.26354e-315
0
14 Logic Display~
6 397 210 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5636 0 0
2
5.90093e-315 0
0
12 IAGO.Nand.4b
94 422 453 0 12 25
0 2 3 4 5 6 7 8 9 10
11 12 13
12 IAGO.Nand.4b
1 0 4752 0
0
2 U1
87 -2 101 6
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
327 0 0
2
45187.7 0
0
66
1 0 2 0 0 4096 0 20 0 0 46 2
382 500
382 601
2 0 3 0 0 4096 0 20 0 0 36 2
410 500
410 574
3 0 4 0 0 4096 0 20 0 0 48 2
445 501
445 546
4 0 5 0 0 4096 0 20 0 0 49 2
481 500
481 522
5 0 6 0 0 4096 0 20 0 0 63 2
369 411
369 315
6 0 7 0 0 4096 0 20 0 0 64 2
387 410
387 302
7 0 8 0 0 4096 0 20 0 0 65 2
405 410
405 287
8 0 9 0 0 4096 0 20 0 0 66 2
422 410
422 274
9 0 10 0 0 4096 0 20 0 0 50 4
450 410
450 392
456 392
456 377
10 0 11 0 0 4096 0 20 0 0 51 4
463 410
463 379
469 379
469 364
11 0 12 0 0 4096 0 20 0 0 52 4
478 410
478 364
484 364
484 349
12 0 13 0 0 4096 0 20 0 0 53 4
489 411
489 351
495 351
495 336
0 0 10 0 0 8448 0 0 0 0 0 5
299 333
339 333
339 380
299 380
299 334
0 0 6 0 0 256 0 0 0 0 0 5
290 269
330 269
330 316
290 316
290 270
1 0 13 0 0 4096 0 1 0 0 53 2
979 447
979 336
2 0 9 0 0 4096 0 1 0 0 17 2
961 447
961 274
0 0 9 0 0 4096 0 0 0 66 0 2
947 274
1219 274
1 0 12 0 0 4096 0 2 0 0 52 2
927 446
927 349
2 0 8 0 0 4096 0 2 0 0 65 2
909 446
909 287
1 0 11 0 0 4096 0 3 0 0 51 2
879 446
879 364
2 0 7 0 0 4096 0 3 0 0 64 2
861 446
861 302
1 0 10 0 0 4096 0 4 0 0 50 2
829 448
829 377
2 0 6 0 0 4096 0 4 0 0 63 2
811 448
811 315
3 0 5 0 0 4096 0 1 0 0 49 2
970 492
970 522
3 0 4 0 0 4096 0 2 0 0 48 2
918 491
918 546
3 0 3 0 0 4096 0 3 0 0 47 2
870 491
870 574
3 0 2 0 0 4096 0 4 0 0 46 2
820 493
820 601
1 0 13 0 0 0 0 5 0 0 53 2
718 228
718 336
1 0 12 0 0 4096 0 6 0 0 52 2
684 227
684 349
1 0 11 0 0 4096 0 7 0 0 51 2
646 228
646 364
1 0 10 0 0 4096 0 8 0 0 50 2
608 228
608 377
4 0 10 0 0 0 0 9 0 0 50 2
548 237
548 377
3 0 11 0 0 0 0 9 0 0 51 2
554 237
554 364
2 0 12 0 0 0 0 9 0 0 52 2
560 237
560 349
1 0 13 0 0 0 0 9 0 0 53 2
566 237
566 336
0 0 3 0 0 4096 0 0 0 47 0 2
639 574
311 574
0 0 14 0 0 8576 0 0 0 0 0 5
1193 514
1260 514
1260 609
1195 609
1195 515
4 0 2 0 0 0 0 14 0 0 46 2
1166 498
1166 601
3 0 3 0 0 0 0 14 0 0 47 2
1172 498
1172 574
2 0 4 0 0 0 0 14 0 0 48 2
1178 498
1178 546
1 0 5 0 0 0 0 14 0 0 49 2
1184 498
1184 522
1 0 2 0 0 4096 0 13 0 0 46 2
1031 479
1031 601
1 0 3 0 0 0 0 12 0 0 47 2
1065 478
1065 574
1 0 4 0 0 4096 0 11 0 0 48 2
1097 477
1097 546
1 0 5 0 0 4096 0 10 0 0 49 2
1128 478
1128 522
0 0 2 0 0 4224 0 0 0 0 0 2
312 601
1222 601
0 0 3 0 0 4224 0 0 0 0 0 2
636 574
1222 574
0 0 4 0 0 4224 0 0 0 0 0 2
311 546
1222 546
0 0 5 0 0 4224 0 0 0 0 0 2
310 522
1222 522
0 0 10 0 0 8320 0 0 0 13 0 3
318 380
318 377
1215 377
0 0 11 0 0 4224 0 0 0 0 0 2
310 364
1215 364
0 0 12 0 0 4224 0 0 0 0 0 2
312 349
1214 349
0 0 13 0 0 4224 0 0 0 0 0 2
310 336
1216 336
0 0 6 0 0 0 0 0 0 63 14 3
318 315
308 315
308 316
4 0 6 0 0 0 0 15 0 0 63 2
341 244
341 315
3 0 7 0 0 0 0 15 0 0 64 2
347 244
347 302
2 0 8 0 0 0 0 15 0 0 65 2
353 244
353 287
1 0 9 0 0 0 0 15 0 0 66 2
359 244
359 274
1 0 6 0 0 0 0 19 0 0 63 2
397 228
397 315
1 0 7 0 0 0 0 18 0 0 64 2
431 227
431 302
1 0 8 0 0 0 0 17 0 0 65 2
463 226
463 287
1 0 9 0 0 0 0 16 0 0 66 2
494 227
494 274
0 0 6 0 0 8320 0 0 0 14 0 3
315 316
315 315
1217 315
0 0 7 0 0 4224 0 0 0 0 0 2
307 302
1218 302
0 0 8 0 0 4224 0 0 0 0 0 2
309 287
1218 287
0 0 9 0 0 4224 0 0 0 0 0 2
307 274
951 274
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1268 544 1321 568
1278 552 1310 568
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
241 273 294 297
251 281 283 297
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1074 399 1135 423
1084 407 1124 423
5 OUT'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
530 127 583 151
540 135 572 151
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
858 217 935 241
868 225 924 241
7 Nand.4b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
240 338 293 362
250 346 282 362
4 BusB
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
