CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
20
11 IAGO.Add.4b
94 924 332 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
11 IAGO.Add.4b
9 0 4224 0
0
2 U7
77 1 91 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3637 0 0
2
45187.8 120
0
13 IAGO.Buffer.4
94 740 333 0 8 17
0 14 15 17 16 10 11 12 13
13 IAGO.Buffer.4
8 0 4224 0
0
2 U6
76 0 90 8
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3226 0 0
2
45187.8 105
0
12 IAGO.Nand.4b
94 543 329 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
12 IAGO.Nand.4b
7 0 4224 0
0
2 U5
87 -2 101 6
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
6966 0 0
2
45187.8 85
0
11 IAGO.Sub.4b
94 361 326 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
11 IAGO.Sub.4b
6 0 4224 0
0
2 U4
80 2 94 10
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
9796 0 0
2
45187.8 15
0
14 Logic Display~
6 909 140 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
45187.8 14
0
14 Logic Display~
6 887 141 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
45187.8 13
0
14 Logic Display~
6 861 140 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
45187.8 12
0
14 Logic Display~
6 839 141 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
45187.8 11
0
8 Hex Key~
166 796 140 0 11 12
0 13 12 11 10 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4681 0 0
2
45187.8 10
0
8 Hex Key~
166 994 146 0 11 12
0 9 8 7 6 0 0 0 0 0
12 67
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9730 0 0
2
45187.8 9
0
14 Logic Display~
6 1122 136 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9874 0 0
2
45187.8 8
0
14 Logic Display~
6 1097 137 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
364 0 0
2
45187.8 7
0
14 Logic Display~
6 1073 137 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3656 0 0
2
45187.8 6
0
14 Logic Display~
6 1051 137 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3131 0 0
2
45187.8 5
0
12 Hex Display~
7 1067 378 0 16 19
10 17 16 15 14 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusU
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6772 0 0
2
45187.8 4
0
14 Logic Display~
6 1189 368 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9557 0 0
2
45187.8 3
0
14 Logic Display~
6 1167 369 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5789 0 0
2
45187.8 2
0
14 Logic Display~
6 1142 369 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7328 0 0
2
45187.8 1
0
14 Logic Display~
6 1117 369 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4799 0 0
2
45187.8 0
0
11 IAGO.ULA.4b
94 199 340 0 1 29
0 0
11 IAGO.ULA.4b
1 0 4224 0
0
2 U8
-82 4 -68 12
0
0
0
0
0
0
29

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
9196 0 0
2
45187.8 0
0
96
14 0 0 0 0 0 0 20 0 0 91 3
243 368
257 368
257 432
13 0 0 0 0 0 0 20 0 0 92 3
256 340
268 340
268 424
9 0 0 0 0 0 0 20 0 0 89 2
188 396
188 451
10 0 0 0 0 0 0 20 0 0 90 2
199 397
199 443
11 0 0 0 0 0 0 20 0 0 91 2
208 396
208 432
12 0 0 0 0 0 0 20 0 0 92 2
218 396
218 424
2 0 0 0 0 0 0 20 0 0 94 2
154 300
154 196
3 0 0 0 0 0 0 20 0 0 95 2
163 302
163 185
4 0 0 0 0 0 0 20 0 0 96 2
172 301
172 177
5 0 0 0 0 0 0 20 0 0 77 2
231 301
231 259
6 0 0 0 0 0 0 20 0 0 78 2
239 300
239 251
7 0 0 0 0 0 0 20 0 0 79 2
248 300
248 240
8 0 0 0 0 0 0 20 0 0 80 2
257 300
257 232
0 0 3 0 0 272 0 0 0 0 0 8
1199 465
1199 416
1243 416
1243 476
1197 476
1197 462
1199 462
1199 461
0 0 4 0 0 272 0 0 0 0 0 5
1195 267
1195 225
1226 225
1226 267
1195 267
0 0 5 0 0 272 0 0 0 0 0 7
1185 159
1185 214
1219 214
1219 156
1186 156
1186 159
1185 159
9 0 6 0 0 16 0 1 0 0 77 2
947 299
947 259
10 0 7 0 0 16 0 1 0 0 78 2
957 298
957 251
11 0 8 0 0 16 0 1 0 0 79 2
965 298
965 240
12 0 9 0 0 16 0 1 0 0 80 2
975 299
975 232
5 0 10 0 0 16 0 1 0 0 93 2
874 299
874 204
6 0 11 0 0 16 0 1 0 0 94 2
884 299
884 196
7 0 12 0 0 16 0 1 0 0 95 2
894 299
894 185
8 0 13 0 0 16 0 1 0 0 96 2
903 299
903 177
5 0 10 0 0 16 0 2 0 0 93 2
695 298
695 204
6 0 11 0 0 16 0 2 0 0 94 2
722 298
722 196
7 0 12 0 0 16 0 2 0 0 95 2
749 300
749 185
8 0 13 0 0 16 0 2 0 0 96 2
778 299
778 177
9 0 6 0 0 16 0 3 0 0 77 2
571 286
571 259
10 0 7 0 0 16 0 3 0 0 78 2
584 286
584 251
11 0 8 0 0 16 0 3 0 0 79 2
599 286
599 240
12 0 9 0 0 16 0 3 0 0 80 2
610 287
610 232
5 0 10 0 0 16 0 3 0 0 93 2
490 287
490 204
6 0 11 0 0 16 0 3 0 0 94 2
508 286
508 196
7 0 12 0 0 16 0 3 0 0 95 2
526 286
526 185
8 0 13 0 0 16 0 3 0 0 96 2
543 286
543 177
9 0 6 0 0 16 0 4 0 0 77 2
388 292
388 259
10 0 7 0 0 16 0 4 0 0 78 2
397 292
397 251
11 0 8 0 0 16 0 4 0 0 79 2
406 291
406 240
12 0 9 0 0 16 0 4 0 0 80 2
416 292
416 232
5 0 10 0 0 16 0 4 0 0 93 2
308 292
308 204
6 0 11 0 0 16 0 4 0 0 94 2
321 293
321 196
7 0 12 0 0 16 0 4 0 0 95 2
334 292
334 185
8 0 13 0 0 16 0 4 0 0 96 2
343 292
343 177
1 0 14 0 0 16 0 1 0 0 89 2
888 377
888 451
2 0 15 0 0 16 0 1 0 0 90 2
915 377
915 443
3 0 16 0 0 16 0 1 0 0 91 2
942 376
942 432
4 0 17 0 0 16 0 1 0 0 92 2
969 376
969 424
1 0 14 0 0 16 0 2 0 0 89 2
695 372
695 451
2 0 15 0 0 16 0 2 0 0 90 2
720 373
720 443
4 0 16 0 0 16 0 2 0 0 91 2
749 372
749 432
3 0 17 0 0 16 0 2 0 0 92 2
777 371
777 424
1 0 14 0 0 16 0 3 0 0 89 2
503 376
503 451
2 0 15 0 0 16 0 3 0 0 90 2
531 376
531 443
3 0 16 0 0 16 0 3 0 0 91 2
566 377
566 432
4 0 17 0 0 16 0 3 0 0 92 2
602 376
602 424
1 0 14 0 0 16 0 4 0 0 89 2
325 372
325 451
2 0 15 0 0 16 0 4 0 0 90 2
352 370
352 443
3 0 16 0 0 16 0 4 0 0 91 2
379 372
379 432
4 0 17 0 0 16 0 4 0 0 92 2
407 371
407 424
4 0 14 0 0 16 0 15 0 0 89 2
1058 402
1058 451
3 0 15 0 0 16 0 15 0 0 90 2
1064 402
1064 443
2 0 16 0 0 16 0 15 0 0 91 2
1070 402
1070 432
1 0 17 0 0 16 0 15 0 0 92 2
1076 402
1076 424
1 0 14 0 0 16 0 19 0 0 89 2
1117 387
1117 451
1 0 15 0 0 16 0 18 0 0 90 2
1142 387
1142 443
1 0 16 0 0 16 0 17 0 0 91 2
1167 387
1167 432
1 0 17 0 0 16 0 16 0 0 92 2
1189 386
1189 424
4 0 6 0 0 16 0 10 0 0 77 2
985 170
985 259
3 0 7 0 0 16 0 10 0 0 78 2
991 170
991 251
2 0 8 0 0 16 0 10 0 0 79 2
997 170
997 240
1 0 9 0 0 16 0 10 0 0 80 2
1003 170
1003 232
1 0 6 0 0 16 0 14 0 0 77 2
1051 155
1051 259
1 0 7 0 0 16 0 13 0 0 78 2
1073 155
1073 251
1 0 8 0 0 16 0 12 0 0 79 2
1097 155
1097 240
1 0 9 0 0 16 0 11 0 0 80 2
1122 154
1122 232
0 0 6 0 0 16 0 0 0 0 0 2
148 259
1204 259
0 0 7 0 0 16 0 0 0 0 0 2
147 251
1205 251
0 0 8 0 0 16 0 0 0 0 0 2
147 240
1203 240
0 0 9 0 0 16 0 0 0 0 0 2
146 232
1204 232
4 0 10 0 0 16 0 9 0 0 93 2
787 164
787 204
3 0 11 0 0 16 0 9 0 0 94 2
793 164
793 196
2 0 12 0 0 16 0 9 0 0 95 2
799 164
799 185
1 0 13 0 0 16 0 9 0 0 96 2
805 164
805 177
1 0 10 0 0 16 0 8 0 0 93 2
839 159
839 204
1 0 11 0 0 16 0 7 0 0 94 2
861 158
861 196
1 0 12 0 0 16 0 6 0 0 95 2
887 159
887 185
1 0 13 0 0 16 0 5 0 0 96 2
909 158
909 177
0 0 14 0 0 16 0 0 0 0 0 2
147 451
1203 451
0 0 15 0 0 16 0 0 0 0 0 2
146 443
1204 443
0 0 16 0 0 16 0 0 0 0 0 2
146 432
1202 432
0 0 17 0 0 16 0 0 0 0 0 2
145 424
1203 424
1 0 10 0 0 16 0 20 0 0 0 3
145 301
145 204
1200 204
0 0 11 0 0 16 0 0 0 0 0 2
143 196
1201 196
0 0 12 0 0 16 0 0 0 0 0 2
143 185
1199 185
0 0 13 0 0 16 0 0 0 0 0 2
142 177
1200 177
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
917 103 970 127
927 111 959 127
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1104 303 1149 327
1114 311 1138 327
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1241 430 1294 454
1251 438 1283 454
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1226 231 1279 255
1236 239 1268 255
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1222 167 1275 191
1232 175 1264 191
4 BusA
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
