CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
11
14 Logic Display~
6 1170 296 0 1 2
10 0
0
0 0 53856 270
6 100MEG
3 -16 45 -8
1 S
-2 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7678 0 0
2
45200.5 0
0
13 IAGO.Decode1b
94 362 347 0 3 7
0 8 7 11
13 IAGO.Decode1b
3 0 4224 0
0
2 U3
77 -9 91 -1
0
0
0
0
0
0
7

0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
961 0 0
2
45200.5 8
0
14 Logic Display~
6 285 135 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
45200.5 7
0
14 Logic Display~
6 279 297 0 1 2
10 11
0
0 0 53856 90
6 100MEG
3 -16 45 -8
1 S
-6 -15 1 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
45200.5 6
0
14 Logic Display~
6 328 132 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
45200.5 5
0
9 2-In AND~
219 664 455 0 3 22
0 8 3 10
0
0 0 96 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8885 0 0
2
45200.5 4
0
9 2-In AND~
219 771 455 0 3 22
0 7 4 9
0
0 0 96 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3780 0 0
2
45200.5 3
0
8 2-In OR~
219 712 512 0 3 22
0 9 10 2
0
0 0 96 270
6 74LS32
-21 -24 21 -16
3 U1A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9265 0 0
2
45200.5 2
0
12 Hex Display~
7 1152 525 0 16 19
10 2 14 15 16 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9442 0 0
2
45200.5 1
0
8 Hex Key~
166 371 143 0 11 12
0 4 3 12 13 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 I0O1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9424 0 0
2
45200.5 0
0
11 IAGO.Mux2x1
94 1010 305 0 1 9
0 0
11 IAGO.Mux2x1
1 0 4224 0
0
2 U4
-90 -6 -76 2
0
0
0
0
0
0
9

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
9968 0 0
2
45200.5 0
0
26
2 0 0 0 0 0 0 11 0 0 25 2
964 265
964 209
3 0 0 0 0 0 0 11 0 0 26 2
1046 265
1046 188
0 1 0 0 0 0 0 0 1 0 0 4
1082 309
1118 309
1118 300
1154 300
1 0 0 0 0 0 0 11 0 0 22 2
1010 339
1010 561
1 0 2 0 0 16 0 9 0 0 22 2
1161 549
1161 561
2 0 3 0 0 16 0 10 0 0 25 2
374 167
374 209
1 0 4 0 0 16 0 10 0 0 26 2
380 167
380 188
0 0 5 0 0 272 0 0 0 0 0 5
1160 369
1160 435
1213 435
1213 369
1160 369
0 0 6 0 0 272 0 0 0 0 0 5
1159 168
1159 225
1213 225
1213 168
1159 168
3 0 2 0 0 16 0 8 0 0 22 2
715 542
715 561
1 0 7 0 0 16 0 7 0 0 24 2
778 433
778 387
2 0 4 0 0 16 0 7 0 0 26 2
760 433
760 188
2 0 3 0 0 16 0 6 0 0 25 2
653 433
653 209
1 0 8 0 0 16 0 6 0 0 23 2
671 433
671 416
3 1 9 0 0 16 0 7 8 0 0 4
769 478
769 491
724 491
724 496
3 2 10 0 0 16 0 6 8 0 0 4
662 478
662 490
706 490
706 496
1 0 8 0 0 16 0 2 0 0 23 2
331 380
331 416
2 0 7 0 0 16 0 2 0 0 24 2
394 381
394 387
1 3 11 0 0 16 0 4 2 0 0 3
294 300
294 303
362 303
1 0 3 0 0 16 0 5 0 0 25 2
328 150
328 209
1 0 4 0 0 16 0 3 0 0 26 2
285 153
285 188
0 0 2 0 0 16 0 0 0 0 0 2
281 561
1171 561
0 0 8 0 0 16 0 0 0 0 0 2
275 416
1174 416
0 0 7 0 0 16 0 0 0 0 0 2
271 387
1175 387
0 0 3 0 0 16 0 0 0 0 0 2
260 209
1175 209
0 0 4 0 0 16 0 0 0 0 0 2
257 188
1176 188
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1171 546 1200 570
1181 554 1189 570
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1175 402 1212 426
1185 410 1201 426
2 M1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1178 371 1215 395
1188 379 1204 395
2 M0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1176 192 1213 216
1186 200 1202 216
2 I1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1177 171 1214 195
1187 179 1203 195
2 I0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
