CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
9961490 0
0
6 Title:
5 Name:
0
0
0
21
14 Logic Display~
6 824 354 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5108 0 0
2
45187.7 0
0
14 Logic Display~
6 804 356 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3320 0 0
2
45187.7 0
0
14 Logic Display~
6 785 357 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
45187.7 0
0
14 Logic Display~
6 765 358 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3557 0 0
2
45187.7 0
0
7 Ground~
168 735 394 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7246 0 0
2
45187.7 0
0
11 IAGO.Add.1b
94 647 381 0 1 11
0 0
11 IAGO.Add.1b
4 0 4224 0
0
2 U4
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3916 0 0
2
45187.7 0
0
11 IAGO.Add.1b
94 477 378 0 1 11
0 0
11 IAGO.Add.1b
3 0 4224 0
0
2 U3
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
614 0 0
2
45187.7 0
0
11 IAGO.Add.1b
94 308 375 0 1 11
0 0
11 IAGO.Add.1b
2 0 4224 0
0
2 U2
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
8494 0 0
2
45187.7 0
0
14 Logic Display~
6 23 355 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Ts3
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
774 0 0
2
45187.7 0
0
8 Hex Key~
166 364 95 0 11 12
0 14 15 16 17 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
715 0 0
2
45187.7 0
0
8 Hex Key~
166 140 98 0 11 12
0 4 3 2 18 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
3281 0 0
2
45187.7 0
0
12 Hex Display~
7 861 372 0 16 19
10 19 20 21 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusW
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3593 0 0
2
45187.7 0
0
14 Logic Display~
6 400 97 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
7233 0 0
2
45187.7 3
0
14 Logic Display~
6 433 96 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3410 0 0
2
45187.7 2
0
14 Logic Display~
6 463 96 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3616 0 0
2
45187.7 1
0
14 Logic Display~
6 495 96 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
5202 0 0
2
45187.7 0
0
14 Logic Display~
6 277 97 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9145 0 0
2
45187.7 0
0
14 Logic Display~
6 245 97 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9815 0 0
2
45187.7 0
0
14 Logic Display~
6 215 97 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4766 0 0
2
45187.7 0
0
14 Logic Display~
6 182 98 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8325 0 0
2
45187.7 0
0
11 IAGO.Add.1b
94 119 372 0 1 11
0 0
11 IAGO.Add.1b
1 0 4224 0
0
2 U1
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
7196 0 0
2
45185.7 0
0
55
1 0 0 0 0 0 0 1 0 0 51 2
824 372
824 442
1 0 0 0 0 0 0 2 0 0 43 2
804 374
804 461
1 0 0 0 0 0 0 3 0 0 42 2
785 375
785 477
1 0 0 0 0 0 0 4 0 0 48 2
765 376
765 496
3 0 0 0 0 0 0 6 0 0 47 2
692 348
692 240
2 0 0 0 0 0 0 6 0 0 55 2
592 348
592 150
5 1 0 0 0 0 0 6 5 0 0 3
715 385
715 388
735 388
1 0 0 0 0 0 0 6 0 0 51 2
647 415
647 442
5 4 0 0 0 0 0 7 6 0 0 3
545 382
545 381
570 381
2 0 0 0 0 0 0 7 0 0 54 2
422 345
422 169
3 0 0 0 0 0 0 7 0 0 46 2
522 345
522 259
1 0 0 0 0 0 0 7 0 0 50 2
477 412
477 461
5 4 0 0 0 0 0 8 7 0 0 3
376 379
376 378
400 378
2 0 0 0 0 0 0 8 0 0 53 2
253 342
253 185
3 0 0 0 0 0 0 8 0 0 45 3
353 342
370 342
370 275
1 0 0 0 0 0 0 8 0 0 49 2
308 409
308 477
5 4 0 0 0 0 0 21 8 0 0 3
187 376
187 375
231 375
1 4 0 0 0 0 0 9 21 0 0 3
23 373
23 372
42 372
1 0 0 0 0 0 0 21 0 0 48 2
119 406
119 496
2 0 0 0 0 0 0 21 0 0 52 2
64 339
64 204
3 0 0 0 0 0 0 21 0 0 44 2
164 339
164 294
4 0 0 0 0 0 0 10 0 0 44 2
355 119
355 294
3 0 0 0 0 0 0 10 0 0 45 2
361 119
361 275
2 0 0 0 0 0 0 10 0 0 46 2
367 119
367 259
1 0 0 0 0 0 0 10 0 0 47 2
373 119
373 240
1 0 0 0 0 0 0 13 0 0 44 2
400 115
400 294
1 0 0 0 0 0 0 14 0 0 45 2
433 114
433 275
1 0 0 0 0 0 0 15 0 0 46 2
463 114
463 259
1 0 0 0 0 0 0 16 0 0 47 2
495 114
495 240
4 0 0 0 0 0 0 12 0 0 48 2
852 396
852 496
3 0 0 0 0 0 0 12 0 0 42 2
858 396
858 477
2 0 0 0 0 0 0 12 0 0 43 2
864 396
864 461
1 0 0 0 0 0 0 12 0 0 51 2
870 396
870 442
4 0 0 0 0 0 0 11 0 0 52 2
131 122
131 204
3 0 0 0 0 0 0 11 0 0 53 2
137 122
137 185
2 0 3 0 0 4096 0 11 0 0 54 2
143 122
143 169
1 0 4 0 0 4096 0 11 0 0 55 2
149 122
149 150
1 0 2 0 0 4096 0 20 0 0 52 2
182 116
182 204
1 0 5 0 0 4096 0 19 0 0 53 2
215 115
215 185
1 0 3 0 0 4096 0 18 0 0 54 2
245 115
245 169
1 0 4 0 0 4096 0 17 0 0 55 2
277 115
277 150
0 0 6 0 0 4096 0 0 0 49 0 2
730 477
897 477
0 0 7 0 0 4096 0 0 0 50 0 2
726 461
898 461
0 0 8 0 0 4224 0 0 0 0 0 2
18 294
727 294
0 0 9 0 0 4224 0 0 0 0 0 2
17 275
729 275
0 0 10 0 0 4224 0 0 0 0 0 2
16 259
725 259
0 0 11 0 0 4224 0 0 0 0 0 2
15 240
727 240
0 0 12 0 0 4224 0 0 0 0 0 2
23 496
897 496
0 0 6 0 0 4224 0 0 0 0 0 2
22 477
734 477
0 0 7 0 0 4224 0 0 0 0 0 2
21 461
730 461
0 0 13 0 0 4224 0 0 0 0 0 2
20 442
899 442
0 0 2 0 0 4224 0 0 0 0 0 2
11 204
720 204
0 0 5 0 0 4224 0 0 0 0 0 2
10 185
722 185
0 0 3 0 0 4224 0 0 0 0 0 2
9 169
718 169
0 0 4 0 0 4224 0 0 0 0 0 2
8 150
720 150
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
788 294 849 318
798 302 838 318
5 OUT's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
273 25 326 49
283 33 315 49
4 IN's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
