CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
15
14 Logic Display~
6 320 159 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5130 0 0
2
45186.5 13
0
14 Logic Display~
6 354 158 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
45186.5 12
0
14 Logic Display~
6 386 157 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
45186.5 11
0
14 Logic Display~
6 417 158 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
45186.5 10
0
14 Logic Display~
6 739 326 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
45186.5 9
0
14 Logic Display~
6 708 325 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
45186.5 8
0
14 Logic Display~
6 676 326 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
45186.5 7
0
14 Logic Display~
6 642 327 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
45186.5 6
0
9 Inverter~
13 427 347 0 2 22
0 5 9
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4747 0 0
2
45186.5 5
0
9 Inverter~
13 457 346 0 2 22
0 6 10
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
972 0 0
2
45186.5 4
0
9 Inverter~
13 488 346 0 2 22
0 7 11
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3472 0 0
2
45186.5 3
0
9 Inverter~
13 519 346 0 2 22
0 8 12
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9998 0 0
2
45186.5 2
0
12 Hex Display~
7 786 340 0 18 19
10 12 11 10 9 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusX
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3536 0 0
2
45186.5 1
0
8 Hex Key~
166 273 169 0 11 12
0 8 7 6 5 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4597 0 0
2
45186.5 0
0
13 IAGO.Buffer.4
94 327 339 0 1 17
0 0
13 IAGO.Buffer.4
1 0 4736 0
0
2 U2
76 0 90 8
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3835 0 0
2
45186.5 0
0
43
1 0 0 0 0 0 0 15 0 0 32 2
282 378
282 467
2 0 0 0 0 0 0 15 0 0 33 2
307 379
307 440
4 0 0 0 0 0 0 15 0 0 34 2
336 378
336 412
3 0 0 0 0 0 0 15 0 0 35 2
364 377
364 388
5 0 0 0 0 0 0 15 0 0 40 2
282 304
282 297
6 0 0 0 0 0 0 15 0 0 41 2
309 304
309 268
7 0 0 0 0 0 0 15 0 0 42 4
336 306
336 259
347 259
347 244
8 0 0 0 0 0 0 15 0 0 43 4
365 305
365 238
376 238
376 223
0 0 2 0 0 272 0 0 0 0 0 5
421 199
563 199
563 494
415 494
415 400
0 0 3 0 0 272 0 0 0 0 0 5
804 380
871 380
871 475
806 475
806 381
0 0 4 0 0 272 0 0 0 0 0 5
190 207
257 207
257 302
192 302
192 208
4 0 5 0 0 16 0 14 0 0 40 2
264 193
264 297
3 0 6 0 0 16 0 14 0 0 41 2
270 193
270 268
2 0 7 0 0 16 0 14 0 0 42 2
276 193
276 244
1 0 8 0 0 16 0 14 0 0 43 2
282 193
282 223
4 0 9 0 0 16 0 13 0 0 32 2
777 364
777 467
3 0 10 0 0 16 0 13 0 0 33 2
783 364
783 440
2 0 11 0 0 16 0 13 0 0 34 2
789 364
789 412
1 0 12 0 0 16 0 13 0 0 35 2
795 364
795 388
2 0 9 0 0 16 0 9 0 0 32 2
430 365
430 467
0 1 5 0 0 16 0 0 9 40 0 3
429 297
430 297
430 329
2 0 10 0 0 16 0 10 0 0 33 2
460 364
460 440
0 1 6 0 0 16 0 0 10 41 0 3
462 268
460 268
460 328
2 0 11 0 0 16 0 11 0 0 34 2
491 364
491 412
0 1 7 0 0 16 0 0 11 42 0 3
489 244
491 244
491 328
2 0 12 0 0 16 0 12 0 0 35 2
522 364
522 388
0 1 8 0 0 16 0 0 12 43 0 3
520 223
522 223
522 328
1 0 9 0 0 16 0 8 0 0 32 2
642 345
642 467
1 0 10 0 0 16 0 7 0 0 33 2
676 344
676 440
1 0 11 0 0 16 0 6 0 0 34 2
708 343
708 412
1 0 12 0 0 16 0 5 0 0 35 2
739 344
739 388
0 0 9 0 0 16 0 0 0 0 0 2
249 467
833 467
0 0 10 0 0 16 0 0 0 0 0 2
247 440
833 440
0 0 11 0 0 16 0 0 0 0 0 2
245 412
833 412
0 0 12 0 0 16 0 0 0 0 0 2
242 388
833 388
1 0 5 0 0 16 0 1 0 0 40 2
320 177
320 297
1 0 6 0 0 16 0 2 0 0 41 2
354 176
354 268
1 0 7 0 0 16 0 3 0 0 42 2
386 175
386 244
1 0 8 0 0 16 0 4 0 0 43 2
417 176
417 223
0 0 5 0 0 16 0 0 0 0 0 2
238 297
591 297
0 0 6 0 0 16 0 0 0 0 0 2
235 268
591 268
0 0 7 0 0 16 0 0 0 0 0 2
232 244
590 244
0 0 8 0 0 16 0 0 0 0 0 2
230 223
592 223
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
456 169 557 193
466 177 546 193
10 Buffer.4b.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
813 351 866 375
823 359 855 375
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
197 179 250 203
207 187 239 203
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
701 261 762 285
711 269 751 285
5 OUT'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
322 94 375 118
332 102 364 118
4 IN'S
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
