CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
19
14 Logic Display~
6 980 263 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5523 0 0
2
45187.8 0
0
14 Logic Display~
6 1005 263 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3330 0 0
2
45187.8 0
0
14 Logic Display~
6 1030 263 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3465 0 0
2
45187.8 0
0
14 Logic Display~
6 1052 262 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 U0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8396 0 0
2
45187.8 0
0
12 Hex Display~
7 930 272 0 16 19
10 14 13 12 11 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusU
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3685 0 0
2
45187.8 0
0
14 Logic Display~
6 914 31 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7849 0 0
2
45187.8 0
0
14 Logic Display~
6 936 31 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6343 0 0
2
45187.8 0
0
14 Logic Display~
6 960 31 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7376 0 0
2
45187.8 0
0
14 Logic Display~
6 985 30 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9156 0 0
2
45187.8 0
0
8 Hex Key~
166 857 40 0 11 12
0 6 5 4 3 0 0 0 0 0
12 67
0
0 0 4656 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
5776 0 0
2
45187.8 0
0
8 Hex Key~
166 659 34 0 11 12
0 10 9 8 7 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7207 0 0
2
45187.8 0
0
14 Logic Display~
6 702 35 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4459 0 0
2
45187.8 0
0
14 Logic Display~
6 724 34 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3760 0 0
2
45187.8 0
0
14 Logic Display~
6 750 35 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
754 0 0
2
45187.8 0
0
14 Logic Display~
6 772 34 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9767 0 0
2
45187.8 0
0
11 IAGO.Sub.4b
94 224 220 0 12 25
0 11 12 13 14 7 8 9 10 3
4 5 6
11 IAGO.Sub.4b
1 0 4240 0
0
2 U4
80 2 94 10
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
7978 0 0
2
45187.7 0
0
12 IAGO.Nand.4b
94 406 223 0 12 25
0 11 12 13 14 7 8 9 10 3
4 5 6
12 IAGO.Nand.4b
2 0 4240 0
0
2 U5
87 -2 101 6
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3142 0 0
2
45187.7 0
0
13 IAGO.Buffer.4
94 603 227 0 8 17
0 11 12 14 13 7 8 9 10
13 IAGO.Buffer.4
3 0 4240 0
0
2 U6
76 0 90 8
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3284 0 0
2
45186.5 0
0
11 IAGO.Add.4b
94 787 226 0 12 25
0 11 12 13 14 7 8 9 10 3
4 5 6
11 IAGO.Add.4b
4 0 4240 0
0
2 U7
77 1 91 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
659 0 0
2
45187.7 0
0
83
0 0 0 0 0 256 0 0 0 0 0 8
1062 359
1062 310
1106 310
1106 370
1060 370
1060 356
1062 356
1062 355
0 0 0 0 0 256 0 0 0 0 0 5
1058 161
1058 119
1089 119
1089 161
1058 161
0 0 0 0 0 256 0 0 0 0 0 7
1048 53
1048 108
1082 108
1082 50
1049 50
1049 53
1048 53
9 0 3 0 0 4096 0 19 0 0 64 2
810 193
810 153
10 0 4 0 0 4096 0 19 0 0 65 2
820 192
820 145
11 0 5 0 0 4096 0 19 0 0 66 2
828 192
828 134
12 0 6 0 0 4096 0 19 0 0 67 2
838 193
838 126
5 0 7 0 0 4096 0 19 0 0 80 2
737 193
737 98
6 0 8 0 0 4096 0 19 0 0 81 2
747 193
747 90
7 0 9 0 0 4096 0 19 0 0 82 2
757 193
757 79
8 0 10 0 0 4096 0 19 0 0 83 2
766 193
766 71
5 0 7 0 0 0 0 18 0 0 80 2
558 192
558 98
6 0 8 0 0 0 0 18 0 0 81 2
585 192
585 90
7 0 9 0 0 4096 0 18 0 0 82 2
612 194
612 79
8 0 10 0 0 0 0 18 0 0 83 2
641 193
641 71
9 0 3 0 0 0 0 17 0 0 64 2
434 180
434 153
10 0 4 0 0 0 0 17 0 0 65 2
447 180
447 145
11 0 5 0 0 0 0 17 0 0 66 2
462 180
462 134
12 0 6 0 0 0 0 17 0 0 67 2
473 181
473 126
5 0 7 0 0 0 0 17 0 0 80 2
353 181
353 98
6 0 8 0 0 0 0 17 0 0 81 2
371 180
371 90
7 0 9 0 0 0 0 17 0 0 82 2
389 180
389 79
8 0 10 0 0 0 0 17 0 0 83 2
406 180
406 71
9 0 3 0 0 0 0 16 0 0 64 2
251 186
251 153
10 0 4 0 0 0 0 16 0 0 65 2
260 186
260 145
11 0 5 0 0 0 0 16 0 0 66 2
269 185
269 134
12 0 6 0 0 0 0 16 0 0 67 2
279 186
279 126
5 0 7 0 0 0 0 16 0 0 80 2
171 186
171 98
6 0 8 0 0 0 0 16 0 0 81 2
184 187
184 90
7 0 9 0 0 0 0 16 0 0 82 2
197 186
197 79
8 0 10 0 0 0 0 16 0 0 83 2
206 186
206 71
1 0 11 0 0 4096 0 19 0 0 76 2
751 271
751 345
2 0 12 0 0 4096 0 19 0 0 77 2
778 271
778 337
3 0 13 0 0 4096 0 19 0 0 78 2
805 270
805 326
4 0 14 0 0 4096 0 19 0 0 79 2
832 270
832 318
1 0 11 0 0 4096 0 18 0 0 76 2
558 266
558 345
2 0 12 0 0 4096 0 18 0 0 77 2
583 267
583 337
4 0 13 0 0 4096 0 18 0 0 78 2
612 266
612 326
3 0 14 0 0 4096 0 18 0 0 79 2
640 265
640 318
1 0 11 0 0 0 0 17 0 0 76 2
366 270
366 345
2 0 12 0 0 0 0 17 0 0 77 2
394 270
394 337
3 0 13 0 0 0 0 17 0 0 78 2
429 271
429 326
4 0 14 0 0 0 0 17 0 0 79 2
465 270
465 318
1 0 11 0 0 0 0 16 0 0 76 2
188 266
188 345
2 0 12 0 0 4096 0 16 0 0 77 2
215 264
215 337
3 0 13 0 0 0 0 16 0 0 78 2
242 266
242 326
4 0 14 0 0 0 0 16 0 0 79 2
270 265
270 318
4 0 11 0 0 0 0 5 0 0 76 2
921 296
921 345
3 0 12 0 0 0 0 5 0 0 77 2
927 296
927 337
2 0 13 0 0 0 0 5 0 0 78 2
933 296
933 326
1 0 14 0 0 0 0 5 0 0 79 2
939 296
939 318
1 0 11 0 0 0 0 1 0 0 76 2
980 281
980 345
1 0 12 0 0 0 0 2 0 0 77 2
1005 281
1005 337
1 0 13 0 0 0 0 3 0 0 78 2
1030 281
1030 326
1 0 14 0 0 0 0 4 0 0 79 2
1052 280
1052 318
4 0 3 0 0 4096 0 10 0 0 64 2
848 64
848 153
3 0 4 0 0 4096 0 10 0 0 65 2
854 64
854 145
2 0 5 0 0 4096 0 10 0 0 66 2
860 64
860 134
1 0 6 0 0 0 0 10 0 0 67 2
866 64
866 126
1 0 3 0 0 4096 0 6 0 0 64 2
914 49
914 153
1 0 4 0 0 4096 0 7 0 0 65 2
936 49
936 145
1 0 5 0 0 4096 0 8 0 0 66 2
960 49
960 134
1 0 6 0 0 4096 0 9 0 0 67 2
985 48
985 126
0 0 3 0 0 4224 0 0 0 0 0 2
11 153
1067 153
0 0 4 0 0 4224 0 0 0 0 0 2
10 145
1068 145
0 0 5 0 0 4224 0 0 0 0 0 2
10 134
1066 134
0 0 6 0 0 4224 0 0 0 0 0 2
9 126
1067 126
4 0 7 0 0 0 0 11 0 0 80 2
650 58
650 98
3 0 8 0 0 0 0 11 0 0 81 2
656 58
656 90
2 0 9 0 0 0 0 11 0 0 82 2
662 58
662 79
1 0 10 0 0 0 0 11 0 0 83 2
668 58
668 71
1 0 7 0 0 0 0 12 0 0 80 2
702 53
702 98
1 0 8 0 0 0 0 13 0 0 81 2
724 52
724 90
1 0 9 0 0 0 0 14 0 0 82 2
750 53
750 79
1 0 10 0 0 0 0 15 0 0 83 2
772 52
772 71
0 0 11 0 0 4224 0 0 0 0 0 2
10 345
1066 345
0 0 12 0 0 4224 0 0 0 0 0 2
9 337
1067 337
0 0 13 0 0 4224 0 0 0 0 0 2
9 326
1065 326
0 0 14 0 0 4224 0 0 0 0 0 2
8 318
1066 318
0 0 7 0 0 4224 0 0 0 0 0 2
7 98
1063 98
0 0 8 0 0 4224 0 0 0 0 0 2
6 90
1064 90
0 0 9 0 0 4224 0 0 0 0 0 2
6 79
1062 79
0 0 10 0 0 4224 0 0 0 0 0 2
5 71
1063 71
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
780 -3 833 21
790 5 822 21
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
967 197 1012 221
977 205 1001 221
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1104 324 1157 348
1114 332 1146 348
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1089 125 1142 149
1099 133 1131 149
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1085 61 1138 85
1095 69 1127 85
4 BusA
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
