CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
15
14 Logic Display~
6 386 122 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.90093e-315 5.41378e-315
0
14 Logic Display~
6 415 121 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.90093e-315 5.4086e-315
0
8 Hex Key~
166 338 123 0 11 12
0 2 9 10 11 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 S1S0
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
5283 0 0
2
5.90093e-315 5.40342e-315
0
12 Hex Display~
7 831 132 0 16 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 N3N0
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6874 0 0
2
5.90093e-315 5.39824e-315
0
14 Logic Display~
6 780 125 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.90093e-315 5.39306e-315
0
14 Logic Display~
6 753 124 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90093e-315 5.38788e-315
0
14 Logic Display~
6 725 124 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.90093e-315 5.37752e-315
0
14 Logic Display~
6 699 125 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.90093e-315 5.36716e-315
0
9 Inverter~
13 455 199 0 2 22
0 9 8
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3751 0 0
2
5.90093e-315 5.3568e-315
0
9 Inverter~
13 482 199 0 2 22
0 2 7
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4292 0 0
2
5.90093e-315 5.34643e-315
0
9 2-In AND~
219 539 269 0 3 22
0 8 7 6
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6118 0 0
2
5.90093e-315 5.32571e-315
0
9 2-In AND~
219 537 318 0 3 22
0 8 2 5
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
34 0 0
2
5.90093e-315 5.30499e-315
0
9 2-In AND~
219 537 372 0 3 22
0 9 7 4
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6357 0 0
2
5.90093e-315 5.26354e-315
0
9 2-In AND~
219 537 422 0 3 22
0 9 2 3
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
319 0 0
2
5.90093e-315 0
0
13 IAGO.Decode.2
94 589 536 0 1 13
0 0
13 IAGO.Decode.2
1 0 4224 0
0
0
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 0 0 0 0
1 U
3976 0 0
2
45187.8 0
0
35
1 0 0 0 0 0 0 15 0 0 33 3
539 578
539 608
699 608
2 0 0 0 0 0 0 15 0 0 32 3
561 579
561 600
725 600
3 0 0 0 0 0 0 15 0 0 31 3
589 580
589 593
753 593
4 0 0 0 0 0 0 15 0 0 30 3
623 579
623 586
780 586
6 0 0 0 0 0 0 15 0 0 34 3
621 489
621 468
415 468
5 0 0 0 0 0 0 15 0 0 35 3
540 488
540 478
386 478
0 0 2 0 0 12672 0 0 0 0 25 5
359 171
359 650
807 650
807 156
356 156
3 0 3 0 0 4096 0 14 0 0 33 2
558 422
699 422
3 0 4 0 0 4096 0 13 0 0 32 2
558 372
725 372
3 0 5 0 0 4096 0 12 0 0 31 2
558 318
753 318
3 0 6 0 0 4096 0 11 0 0 30 2
560 269
780 269
2 0 7 0 0 4352 0 13 0 0 16 2
513 381
485 381
2 0 7 0 0 4352 0 11 0 0 16 2
515 278
485 278
1 0 8 0 0 4352 0 11 0 0 17 2
515 260
458 260
1 0 8 0 0 0 0 12 0 0 17 2
513 309
458 309
2 0 7 0 0 4480 0 10 0 0 0 2
485 217
485 623
2 0 8 0 0 4480 0 9 0 0 0 2
458 217
458 621
2 0 2 0 0 0 0 12 0 0 34 2
513 327
415 327
1 0 9 0 0 4096 0 13 0 0 35 2
513 363
386 363
2 0 2 0 0 0 0 14 0 0 34 2
513 431
415 431
1 0 9 0 0 0 0 14 0 0 35 2
513 413
386 413
0 1 2 0 0 0 0 0 10 34 0 3
415 143
485 143
485 181
0 1 9 0 0 0 0 0 9 35 0 3
386 150
458 150
458 181
2 0 9 0 0 0 0 3 0 0 35 3
341 147
341 163
386 163
1 0 2 0 0 0 0 3 0 0 34 3
347 147
347 156
415 156
1 0 6 0 0 0 0 4 0 0 30 3
840 156
840 194
780 194
2 0 5 0 0 0 0 4 0 0 31 3
834 156
834 184
753 184
3 0 4 0 0 0 0 4 0 0 32 3
828 156
828 176
725 176
4 0 3 0 0 0 0 4 0 0 33 3
822 156
822 170
699 170
1 0 6 0 0 4224 0 5 0 0 0 2
780 143
780 624
1 0 5 0 0 4224 0 6 0 0 0 2
753 142
753 625
1 0 4 0 0 4224 0 7 0 0 0 2
725 142
725 627
1 0 3 0 0 4224 0 8 0 0 0 2
699 143
699 627
1 0 2 0 0 0 0 2 0 0 0 2
415 139
415 626
1 0 9 0 0 4224 0 1 0 0 0 2
386 140
386 627
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
549 130 642 154
559 138 631 154
9 Decode.2b
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
