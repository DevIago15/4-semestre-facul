CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
-1424 28 -2 779
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
-1256 124 -1143 221
9961490 0
0
6 Title:
5 Name:
0
0
0
19
8 2-In OR~
219 596 392 0 3 22
0 4 3 2
0
0 0 96 0
4 4071
-15 -24 13 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 96293112
65 0 0 0 4 1 2 0
1 U
5130 0 0
2
5.90093e-315 0
0
9 2-In AND~
219 549 474 0 3 22
0 9 8 3
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
391 0 0
2
5.90093e-315 0
0
9 2-In AND~
219 547 423 0 3 22
0 10 7 18
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
3124 0 0
2
5.90093e-315 0
0
9 2-In AND~
219 548 369 0 3 22
0 11 6 19
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 1 0
1 U
3421 0 0
2
5.90093e-315 0
0
9 2-In AND~
219 545 319 0 3 22
0 12 5 4
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8157 0 0
2
5.90093e-315 0
0
12 Hex Display~
7 690 86 0 16 19
10 2 20 21 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
5572 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 639 78 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 358 76 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 327 77 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 288 93 0 11 12
0 14 13 23 24 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 S1S0
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
972 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 55 462 0 11 12
0 8 25 26 27 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3472 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 54 361 0 11 12
0 7 28 29 30 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9998 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 56 260 0 11 12
0 6 31 32 33 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3536 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 53 174 0 11 12
0 5 34 35 36 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I0
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
4597 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 189 87 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 137 88 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 163 87 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 108 88 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90093e-315 0
0
13 IAGO.Decode.2
94 451 219 0 6 13
0 9 10 11 12 13 14
13 IAGO.Decode.2
1 0 4736 0
0
2 U1
74 -5 88 3
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
1 U
317 0 0
2
5.90093e-315 0
0
29
3 0 0 0 0 0 0 3 0 0 0 4
568 423
578 423
578 397
589 397
3 0 0 0 0 0 0 4 0 0 0 4
569 369
577 369
577 389
590 389
1 0 2 0 0 8192 0 6 0 0 25 3
699 110
699 129
639 129
3 2 3 0 0 8320 0 2 1 0 0 3
570 474
583 474
583 401
3 1 4 0 0 8320 0 5 1 0 0 3
566 319
583 319
583 383
3 0 2 0 0 0 0 1 0 0 25 2
629 392
639 392
2 0 5 0 0 4096 0 5 0 0 26 2
521 328
189 328
2 0 6 0 0 4096 0 4 0 0 27 2
524 378
163 378
2 0 7 0 0 4096 0 3 0 0 28 2
523 432
137 432
2 0 8 0 0 4096 0 2 0 0 29 2
525 483
108 483
1 1 9 0 0 4224 0 19 2 0 0 3
401 261
401 465
525 465
2 1 10 0 0 4224 0 19 3 0 0 3
423 262
423 414
523 414
3 1 11 0 0 4224 0 19 4 0 0 3
451 263
451 360
524 360
4 1 12 0 0 4224 0 19 5 0 0 3
485 262
485 310
521 310
0 5 13 0 0 4352 0 0 19 20 0 3
327 164
402 164
402 171
0 6 14 0 0 4352 0 0 19 19 0 3
358 141
483 141
483 172
2 0 13 0 0 256 0 10 0 0 20 3
291 117
291 153
327 153
1 0 14 0 0 256 0 10 0 0 19 3
297 117
297 133
358 133
1 0 14 0 0 4480 0 8 0 0 0 2
358 94
358 645
1 0 13 0 0 4480 0 9 0 0 0 2
327 95
327 644
1 0 8 0 0 0 0 11 0 0 29 3
64 486
64 499
108 499
1 0 7 0 0 0 0 12 0 0 28 3
63 385
63 404
137 404
1 0 6 0 0 0 0 13 0 0 27 3
65 284
65 291
163 291
1 0 5 0 0 0 0 14 0 0 26 3
62 198
62 208
189 208
1 0 2 0 0 4224 0 7 0 0 0 2
639 96
639 643
1 0 5 0 0 4224 0 15 0 0 0 2
189 105
189 644
1 0 6 0 0 4224 0 17 0 0 0 2
163 105
163 645
1 0 7 0 0 4224 0 16 0 0 0 2
137 106
137 647
1 0 8 0 0 4224 0 18 0 0 0 2
108 106
108 647
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
125 21 178 45
135 29 167 45
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
261 20 314 44
271 28 303 44
4 Ctrl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
618 20 663 44
628 28 652 44
3 Out
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
