CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2096 80 3518 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
2264 176 2377 273
42991634 0
0
6 Title:
5 Name:
0
0
0
19
9 2-In AND~
219 972 434 0 3 22
0 4 5 10
0
0 0 112 270
6 74LS08
-21 -24 21 -16
2 A1
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5130 0 0
2
5.90093e-315 5.32571e-315
0
9 2-In AND~
219 920 433 0 3 22
0 6 7 11
0
0 0 112 270
6 74LS08
-21 -24 21 -16
2 A2
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
391 0 0
2
5.90093e-315 5.30499e-315
0
9 2-In AND~
219 872 433 0 3 22
0 8 9 12
0
0 0 112 270
6 74LS08
-21 -24 21 -16
2 A3
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3124 0 0
2
5.90093e-315 5.26354e-315
0
9 2-In AND~
219 822 435 0 3 22
0 2 3 13
0
0 0 112 270
6 74LS08
-21 -24 21 -16
2 A4
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3421 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 718 175 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 684 174 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 646 175 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 608 175 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90093e-315 0
0
8 Hex Key~
166 557 178 0 11 12
0 4 6 8 2 0 0 0 0 0
14 69
0
0 0 4656 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4747 0 0
2
5.90093e-315 0
0
14 Logic Display~
6 1128 425 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90093e-315 5.38788e-315
0
14 Logic Display~
6 1097 424 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90093e-315 5.37752e-315
0
14 Logic Display~
6 1065 425 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90093e-315 5.36716e-315
0
14 Logic Display~
6 1031 426 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90093e-315 5.3568e-315
0
12 Hex Display~
7 1175 439 0 18 19
10 10 11 12 13 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusY
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4597 0 0
2
5.90093e-315 5.34643e-315
0
8 Hex Key~
166 350 185 0 11 12
0 5 7 9 3 0 0 0 0 0
10 65
0
0 0 4656 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3835 0 0
2
5.90093e-315 5.41378e-315
0
14 Logic Display~
6 494 174 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90093e-315 5.32571e-315
0
14 Logic Display~
6 463 173 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90093e-315 5.30499e-315
0
14 Logic Display~
6 431 174 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90093e-315 5.26354e-315
0
14 Logic Display~
6 397 175 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90093e-315 0
0
54
0 0 2 0 0 8464 0 0 0 0 0 5
299 298
339 298
339 345
299 345
299 299
0 0 3 0 0 8448 0 0 0 0 0 5
290 234
330 234
330 281
290 281
290 235
1 0 4 0 0 4096 0 1 0 0 41 2
979 412
979 301
2 0 5 0 0 4096 0 1 0 0 5 2
961 412
961 239
0 0 5 0 0 4096 0 0 0 54 0 2
947 239
1219 239
1 0 6 0 0 4096 0 2 0 0 40 2
927 411
927 314
2 0 7 0 0 4096 0 2 0 0 53 2
909 411
909 252
1 0 8 0 0 4096 0 3 0 0 39 2
879 411
879 329
2 0 9 0 0 4096 0 3 0 0 52 2
861 411
861 267
1 0 2 0 0 4096 0 4 0 0 38 2
829 413
829 342
2 0 3 0 0 4096 0 4 0 0 51 2
811 413
811 280
3 0 10 0 0 4096 0 1 0 0 37 2
970 457
970 487
3 0 11 0 0 4096 0 2 0 0 36 2
918 456
918 511
3 0 12 0 0 4096 0 3 0 0 35 2
870 456
870 539
3 0 13 0 0 4096 0 4 0 0 34 2
820 458
820 566
1 0 4 0 0 0 0 5 0 0 41 2
718 193
718 301
1 0 6 0 0 4096 0 6 0 0 40 2
684 192
684 314
1 0 8 0 0 4096 0 7 0 0 39 2
646 193
646 329
1 0 2 0 0 4096 0 8 0 0 38 2
608 193
608 342
4 0 2 0 0 0 0 9 0 0 38 2
548 202
548 342
3 0 8 0 0 0 0 9 0 0 39 2
554 202
554 329
2 0 6 0 0 0 0 9 0 0 40 2
560 202
560 314
1 0 4 0 0 0 0 9 0 0 41 2
566 202
566 301
0 0 12 0 0 4096 0 0 0 35 0 2
639 539
311 539
0 0 14 0 0 8576 0 0 0 0 0 5
1193 479
1260 479
1260 574
1195 574
1195 480
4 0 13 0 0 0 0 14 0 0 34 2
1166 463
1166 566
3 0 12 0 0 0 0 14 0 0 35 2
1172 463
1172 539
2 0 11 0 0 0 0 14 0 0 36 2
1178 463
1178 511
1 0 10 0 0 0 0 14 0 0 37 2
1184 463
1184 487
1 0 13 0 0 4096 0 13 0 0 34 2
1031 444
1031 566
1 0 12 0 0 0 0 12 0 0 35 2
1065 443
1065 539
1 0 11 0 0 4096 0 11 0 0 36 2
1097 442
1097 511
1 0 10 0 0 4096 0 10 0 0 37 2
1128 443
1128 487
0 0 13 0 0 4224 0 0 0 0 0 2
312 566
1222 566
0 0 12 0 0 4224 0 0 0 0 0 2
636 539
1222 539
0 0 11 0 0 4224 0 0 0 0 0 2
311 511
1222 511
0 0 10 0 0 4224 0 0 0 0 0 2
310 487
1222 487
0 0 2 0 0 8320 0 0 0 1 0 3
318 345
318 342
1215 342
0 0 8 0 0 4224 0 0 0 0 0 2
310 329
1215 329
0 0 6 0 0 4224 0 0 0 0 0 2
312 314
1214 314
0 0 4 0 0 4224 0 0 0 0 0 2
310 301
1216 301
0 0 3 0 0 0 0 0 0 51 2 3
318 280
308 280
308 281
4 0 3 0 0 0 0 15 0 0 51 2
341 209
341 280
3 0 9 0 0 0 0 15 0 0 52 2
347 209
347 267
2 0 7 0 0 0 0 15 0 0 53 2
353 209
353 252
1 0 5 0 0 0 0 15 0 0 54 2
359 209
359 239
1 0 3 0 0 0 0 19 0 0 51 2
397 193
397 280
1 0 9 0 0 0 0 18 0 0 52 2
431 192
431 267
1 0 7 0 0 0 0 17 0 0 53 2
463 191
463 252
1 0 5 0 0 0 0 16 0 0 54 2
494 192
494 239
0 0 3 0 0 8320 0 0 0 2 0 3
315 281
315 280
1217 280
0 0 9 0 0 4224 0 0 0 0 0 2
307 267
1218 267
0 0 7 0 0 4224 0 0 0 0 0 2
309 252
1218 252
0 0 5 0 0 4224 0 0 0 0 0 2
307 239
951 239
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
241 238 294 262
251 246 283 262
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1074 364 1135 388
1084 372 1124 388
5 OUT'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
530 92 583 116
540 100 572 116
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
738 179 815 203
748 187 804 203
7 Nand.4b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
240 303 293 327
250 311 282 327
4 BusB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
