CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 160 30 100 10
-1424 28 -2 779
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
-1256 124 -1143 221
9961490 0
0
6 Title:
5 Name:
0
0
0
27
14 Logic Display~
6 1110 758 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
45190.7 328
0
14 Logic Display~
6 1089 759 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
45190.7 327
0
8 Hex Key~
166 1062 751 0 11 12
0 4 3 221 222 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 Ctrl
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3221 0 0
2
45190.7 326
0
12 IAGO.Mux.4x1
94 880 756 0 7 15
0 4 3 10 11 13 12 5
12 IAGO.Mux.4x1
17 0 4224 0
0
3 U11
68 3 89 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3215 0 0
2
45190.7 292
0
12 IAGO.Mux.4x1
94 699 755 0 7 15
0 4 3 15 14 16 9 6
12 IAGO.Mux.4x1
16 0 4224 0
0
3 U10
68 3 89 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7903 0 0
2
45190.7 258
0
12 IAGO.Mux.4x1
94 505 755 0 7 15
0 4 3 17 18 19 9 7
12 IAGO.Mux.4x1
15 0 4224 0
0
2 U9
71 3 85 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7121 0 0
2
45190.7 224
0
12 Hex Display~
7 1155 797 0 16 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 BusU
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4484 0 0
2
45190.7 223
0
14 Logic Display~
6 1277 787 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
45190.7 222
0
14 Logic Display~
6 1255 788 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
45190.7 221
0
14 Logic Display~
6 1230 788 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
45190.7 220
0
14 Logic Display~
6 1205 788 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
45190.7 219
0
14 Logic Display~
6 1123 55 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
45190.7 218
0
14 Logic Display~
6 1145 55 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
45190.7 217
0
14 Logic Display~
6 1169 55 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
45190.7 216
0
14 Logic Display~
6 1194 54 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
45190.7 215
0
8 Hex Key~
166 1066 64 0 11 12
0 35 34 33 32 0 0 0 0 0
12 67
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6343 0 0
2
45190.7 214
0
8 Hex Key~
166 868 58 0 11 12
0 39 38 37 36 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7376 0 0
2
45190.7 213
0
14 Logic Display~
6 911 59 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
45190.7 212
0
14 Logic Display~
6 933 58 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
45190.7 211
0
14 Logic Display~
6 959 59 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
45190.7 210
0
14 Logic Display~
6 981 58 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
45190.7 209
0
11 IAGO.Sub.4b
94 433 244 0 12 25
0 20 17 15 10 36 37 38 39 32
33 34 35
11 IAGO.Sub.4b
14 0 4224 0
0
2 U4
80 2 94 10
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3760 0 0
2
45190.7 139
0
12 IAGO.Nand.4b
94 615 247 0 12 25
0 21 14 18 11 36 37 38 39 32
33 34 35
12 IAGO.Nand.4b
13 0 4224 0
0
2 U5
87 -2 101 6
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
754 0 0
2
45190.7 119
0
13 IAGO.Buffer.4
94 812 251 0 8 17
0 22 24 12 9 36 37 38 39
13 IAGO.Buffer.4
12 0 4224 0
0
2 U6
76 0 90 8
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
9767 0 0
2
45190.7 104
0
11 IAGO.Add.4b
94 996 250 0 12 25
0 23 19 16 13 36 37 38 39 32
33 34 35
11 IAGO.Add.4b
11 0 4224 0
0
2 U7
77 1 91 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7978 0 0
2
45190.7 34
0
12 IAGO.Mux.4x1
94 320 753 0 7 15
0 4 3 20 21 23 22 8
12 IAGO.Mux.4x1
10 0 4224 0
0
2 U8
71 3 85 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3142 0 0
2
45190.7 0
0
11 IAGO.ULA.4b
94 77 624 0 1 29
0 0
11 IAGO.ULA.4b
1 0 4224 0
0
3 U12
-88 2 -67 10
0
0
0
0
0
0
29

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3284 0 0
2
45190.7 0
0
142
1 0 0 0 0 0 0 27 0 0 69 2
60 681
60 870
2 0 0 0 0 0 0 27 0 0 7 2
68 680
68 862
3 0 0 0 0 0 0 27 0 0 71 2
77 679
77 851
4 0 0 0 0 0 0 27 0 0 72 2
87 681
87 843
14 0 0 0 0 256 0 27 0 0 0 4
116 646
151 646
151 832
257 832
13 0 0 0 0 256 0 27 0 0 23 4
129 624
165 624
165 818
275 818
0 0 0 0 0 0 0 0 0 70 0 2
237 862
21 862
2 0 3 0 0 272 0 4 0 0 22 3
802 778
791 778
791 829
1 0 4 0 0 272 0 4 0 0 23 3
802 756
787 756
787 818
2 0 3 0 0 272 0 5 0 0 22 3
621 777
609 777
609 829
1 0 4 0 0 272 0 5 0 0 23 3
621 755
602 755
602 818
2 0 3 0 0 272 0 6 0 0 22 3
427 777
420 777
420 829
1 0 4 0 0 272 0 6 0 0 23 3
427 755
414 755
414 818
7 0 5 0 0 16 0 4 0 0 72 2
880 800
880 843
7 0 6 0 0 16 0 5 0 0 71 2
699 799
699 851
7 0 7 0 0 16 0 6 0 0 70 2
505 799
505 862
7 0 8 0 0 16 0 26 0 0 69 2
320 797
320 870
2 0 3 0 0 16 0 3 0 0 22 2
1065 775
1065 829
1 0 4 0 0 16 0 3 0 0 23 2
1071 775
1071 818
1 0 3 0 0 272 0 2 0 0 22 2
1089 777
1089 829
1 0 4 0 0 272 0 1 0 0 23 2
1110 776
1110 818
2 0 3 0 0 272 0 26 0 0 0 4
242 775
237 775
237 829
1123 829
1 0 4 0 0 272 0 26 0 0 0 4
242 753
234 753
234 818
1123 818
6 0 9 0 0 16 0 5 0 0 83 2
706 725
706 504
3 0 10 0 0 16 0 4 0 0 76 2
829 725
829 641
4 0 11 0 0 16 0 4 0 0 80 2
860 727
860 566
6 0 12 0 0 16 0 4 0 0 84 2
887 726
887 487
5 0 13 0 0 16 0 4 0 0 88 2
913 726
913 417
4 0 14 0 0 16 0 5 0 0 78 2
679 726
679 595
3 0 15 0 0 16 0 5 0 0 75 2
648 724
648 658
5 0 16 0 0 16 0 5 0 0 87 2
732 725
732 434
3 0 17 0 0 16 0 6 0 0 74 2
454 724
454 670
4 0 18 0 0 16 0 6 0 0 79 2
485 726
485 583
6 0 9 0 0 16 0 6 0 0 83 2
512 725
512 504
5 0 19 0 0 16 0 6 0 0 86 2
538 725
538 446
3 0 20 0 0 16 0 26 0 0 73 2
269 722
269 683
4 0 21 0 0 16 0 26 0 0 77 2
300 724
300 608
6 0 22 0 0 16 0 26 0 0 81 2
327 723
327 529
5 0 23 0 0 16 0 26 0 0 85 2
353 723
353 459
1 0 20 0 0 16 0 22 0 0 73 2
397 290
397 683
2 0 17 0 0 16 0 22 0 0 74 2
424 288
424 670
3 0 15 0 0 16 0 22 0 0 75 2
451 290
451 658
4 0 10 0 0 16 0 22 0 0 76 2
479 289
479 641
1 0 21 0 0 16 0 23 0 0 77 2
575 294
575 608
2 0 14 0 0 16 0 23 0 0 78 2
603 294
603 595
3 0 18 0 0 16 0 23 0 0 79 2
638 295
638 583
4 0 11 0 0 16 0 23 0 0 80 2
674 294
674 566
1 0 22 0 0 16 0 24 0 0 81 2
767 290
767 529
2 0 24 0 0 16 0 24 0 0 82 2
792 291
792 516
4 0 9 0 0 16 0 24 0 0 83 2
821 290
821 504
3 0 12 0 0 16 0 24 0 0 84 2
849 289
849 487
1 0 23 0 0 16 0 25 0 0 85 2
960 295
960 459
2 0 19 0 0 16 0 25 0 0 86 2
987 295
987 446
3 0 16 0 0 16 0 25 0 0 87 2
1014 294
1014 434
4 0 13 0 0 16 0 25 0 0 88 2
1041 294
1041 417
0 0 25 0 0 272 0 0 0 0 0 5
1226 631
1226 694
1294 694
1294 631
1226 631
0 0 26 0 0 272 0 0 0 0 0 5
1226 559
1226 620
1293 620
1293 559
1226 559
0 0 27 0 0 272 0 0 0 0 0 5
1224 543
1224 481
1293 481
1293 547
1224 547
0 0 28 0 0 272 0 0 0 0 0 5
1220 380
1220 472
1291 472
1291 380
1220 380
0 0 29 0 0 272 0 0 0 0 0 8
1287 884
1287 835
1331 835
1331 895
1285 895
1285 881
1287 881
1287 880
4 0 8 0 0 16 0 7 0 0 69 2
1146 821
1146 870
3 0 7 0 0 16 0 7 0 0 70 2
1152 821
1152 862
2 0 6 0 0 16 0 7 0 0 71 2
1158 821
1158 851
1 0 5 0 0 16 0 7 0 0 72 2
1164 821
1164 843
1 0 8 0 0 16 0 11 0 0 69 2
1205 806
1205 870
1 0 7 0 0 16 0 10 0 0 70 2
1230 806
1230 862
1 0 6 0 0 16 0 9 0 0 71 2
1255 806
1255 851
1 0 5 0 0 16 0 8 0 0 72 2
1277 805
1277 843
0 0 8 0 0 16 0 0 0 0 0 2
20 870
1291 870
0 0 7 0 0 16 0 0 0 0 0 2
234 862
1292 862
0 0 6 0 0 16 0 0 0 0 0 2
21 851
1290 851
0 0 5 0 0 16 0 0 0 0 0 2
22 843
1291 843
0 0 20 0 0 16 0 0 0 0 0 2
229 683
1271 683
0 0 17 0 0 16 0 0 0 0 0 2
226 670
1272 670
0 0 15 0 0 16 0 0 0 0 0 2
225 658
1272 658
0 0 10 0 0 16 0 0 0 0 0 2
225 641
1273 641
0 0 21 0 0 16 0 0 0 0 0 2
227 608
1269 608
0 0 14 0 0 16 0 0 0 0 0 2
224 595
1270 595
0 0 18 0 0 16 0 0 0 0 0 2
223 583
1270 583
0 0 11 0 0 16 0 0 0 0 0 2
223 566
1271 566
0 0 22 0 0 16 0 0 0 0 0 2
226 529
1268 529
0 0 24 0 0 16 0 0 0 0 0 2
223 516
1269 516
0 0 9 0 0 16 0 0 0 0 0 2
222 504
1269 504
0 0 12 0 0 16 0 0 0 0 0 2
222 487
1270 487
0 0 23 0 0 16 0 0 0 0 0 2
227 459
1269 459
0 0 19 0 0 16 0 0 0 0 0 2
224 446
1270 446
0 0 16 0 0 16 0 0 0 0 0 2
223 434
1270 434
0 0 13 0 0 16 0 0 0 0 0 2
223 417
1271 417
0 0 30 0 0 272 0 0 0 0 0 5
1267 185
1267 143
1298 143
1298 185
1267 185
0 0 31 0 0 272 0 0 0 0 0 7
1257 77
1257 132
1291 132
1291 74
1258 74
1258 77
1257 77
9 0 32 0 0 16 0 25 0 0 127 2
1019 217
1019 177
10 0 33 0 0 16 0 25 0 0 128 2
1029 216
1029 169
11 0 34 0 0 16 0 25 0 0 129 2
1037 216
1037 158
12 0 35 0 0 16 0 25 0 0 130 2
1047 217
1047 150
5 0 36 0 0 16 0 25 0 0 139 2
946 217
946 122
6 0 37 0 0 16 0 25 0 0 140 2
956 217
956 114
7 0 38 0 0 16 0 25 0 0 141 2
966 217
966 103
8 0 39 0 0 16 0 25 0 0 142 2
975 217
975 95
5 0 36 0 0 16 0 24 0 0 139 2
767 216
767 122
6 0 37 0 0 16 0 24 0 0 140 2
794 216
794 114
7 0 38 0 0 16 0 24 0 0 141 2
821 218
821 103
8 0 39 0 0 16 0 24 0 0 142 2
850 217
850 95
9 0 32 0 0 16 0 23 0 0 127 2
643 204
643 177
10 0 33 0 0 16 0 23 0 0 128 2
656 204
656 169
11 0 34 0 0 16 0 23 0 0 129 2
671 204
671 158
12 0 35 0 0 16 0 23 0 0 130 2
682 205
682 150
5 0 36 0 0 16 0 23 0 0 139 2
562 205
562 122
6 0 37 0 0 16 0 23 0 0 140 2
580 204
580 114
7 0 38 0 0 16 0 23 0 0 141 2
598 204
598 103
8 0 39 0 0 16 0 23 0 0 142 2
615 204
615 95
9 0 32 0 0 16 0 22 0 0 127 2
460 210
460 177
10 0 33 0 0 16 0 22 0 0 128 2
469 210
469 169
11 0 34 0 0 16 0 22 0 0 129 2
478 209
478 158
12 0 35 0 0 16 0 22 0 0 130 2
488 210
488 150
5 0 36 0 0 16 0 22 0 0 139 2
380 210
380 122
6 0 37 0 0 16 0 22 0 0 140 2
393 211
393 114
7 0 38 0 0 16 0 22 0 0 141 2
406 210
406 103
8 0 39 0 0 16 0 22 0 0 142 2
415 210
415 95
4 0 32 0 0 16 0 16 0 0 127 2
1057 88
1057 177
3 0 33 0 0 16 0 16 0 0 128 2
1063 88
1063 169
2 0 34 0 0 16 0 16 0 0 129 2
1069 88
1069 158
1 0 35 0 0 16 0 16 0 0 130 2
1075 88
1075 150
1 0 32 0 0 16 0 12 0 0 127 2
1123 73
1123 177
1 0 33 0 0 16 0 13 0 0 128 2
1145 73
1145 169
1 0 34 0 0 16 0 14 0 0 129 2
1169 73
1169 158
1 0 35 0 0 16 0 15 0 0 130 2
1194 72
1194 150
0 0 32 0 0 16 0 0 0 0 0 2
220 177
1276 177
0 0 33 0 0 16 0 0 0 0 0 2
219 169
1277 169
0 0 34 0 0 16 0 0 0 0 0 2
219 158
1275 158
0 0 35 0 0 16 0 0 0 0 0 2
218 150
1276 150
4 0 36 0 0 16 0 17 0 0 139 2
859 82
859 122
3 0 37 0 0 16 0 17 0 0 140 2
865 82
865 114
2 0 38 0 0 16 0 17 0 0 141 2
871 82
871 103
1 0 39 0 0 16 0 17 0 0 142 2
877 82
877 95
1 0 36 0 0 16 0 18 0 0 139 2
911 77
911 122
1 0 37 0 0 16 0 19 0 0 140 2
933 76
933 114
1 0 38 0 0 16 0 20 0 0 141 2
959 77
959 103
1 0 39 0 0 16 0 21 0 0 142 2
981 76
981 95
0 0 36 0 0 16 0 0 0 0 0 2
216 122
1272 122
0 0 37 0 0 16 0 0 0 0 0 2
215 114
1273 114
0 0 38 0 0 16 0 0 0 0 0 2
215 103
1271 103
0 0 39 0 0 16 0 0 0 0 0 2
214 95
1272 95
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
989 21 1042 45
999 29 1031 45
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1298 149 1351 173
1308 157 1340 173
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1294 85 1347 109
1304 93 1336 109
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1329 849 1382 873
1339 857 1371 873
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1207 731 1252 755
1217 739 1241 755
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1310 643 1363 667
1320 651 1352 667
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1315 660 1360 684
1325 668 1349 684
3 Sub
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1306 559 1359 583
1316 567 1348 583
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1307 575 1360 599
1317 583 1349 599
4 Nand
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1305 480 1358 504
1315 488 1347 504
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1299 497 1368 521
1309 505 1357 521
6 Buffer
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1307 406 1360 430
1317 414 1349 430
4 BusW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1309 424 1354 448
1319 432 1343 448
3 Add
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1041 689 1118 713
1051 697 1107 713
7 Fun��es
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
