CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
8 Hex Key~
166 178 62 0 11 12
0 4 3 12 13 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 I0O1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
972 0 0
2
45200.5 0
0
12 Hex Display~
7 959 444 0 16 19
10 2 14 15 16 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3472 0 0
2
45200.5 0
0
8 2-In OR~
219 519 431 0 3 22
0 9 10 2
0
0 0 112 270
6 74LS32
-21 -24 21 -16
3 U3A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9998 0 0
2
45200.5 0
0
9 2-In AND~
219 578 374 0 3 22
0 7 4 9
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3536 0 0
2
45200.5 0
0
9 2-In AND~
219 471 374 0 3 22
0 8 3 10
0
0 0 112 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4597 0 0
2
45200.5 0
0
14 Logic Display~
6 135 51 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
45200.5 0
0
14 Logic Display~
6 86 216 0 1 2
10 11
0
0 0 53856 90
6 100MEG
3 -16 45 -8
1 S
-6 -15 1 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45200.5 0
0
14 Logic Display~
6 92 54 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 I0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45200.5 0
0
13 IAGO.Decode1b
94 169 266 0 3 7
0 8 7 11
13 IAGO.Decode1b
1 0 4240 0
0
2 U1
77 -9 91 -1
0
0
0
0
0
0
7

0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
9323 0 0
2
45199.7 0
0
22
1 0 2 0 0 4096 0 2 0 0 18 2
968 468
968 480
2 0 3 0 0 4096 0 1 0 0 21 2
181 86
181 128
1 0 4 0 0 4096 0 1 0 0 22 2
187 86
187 107
0 0 5 0 0 4480 0 0 0 0 0 5
967 288
967 354
1020 354
1020 288
967 288
0 0 6 0 0 4480 0 0 0 0 0 5
966 87
966 144
1020 144
1020 87
966 87
3 0 2 0 0 4096 0 3 0 0 18 2
522 461
522 480
1 0 7 0 0 4096 0 4 0 0 20 2
585 352
585 306
2 0 4 0 0 4096 0 4 0 0 22 2
567 352
567 107
2 0 3 0 0 4096 0 5 0 0 21 2
460 352
460 128
1 0 8 0 0 4096 0 5 0 0 19 2
478 352
478 335
3 1 9 0 0 8320 0 4 3 0 0 4
576 397
576 410
531 410
531 415
3 2 10 0 0 8320 0 5 3 0 0 4
469 397
469 409
513 409
513 415
1 0 8 0 0 4096 0 9 0 0 19 2
138 299
138 335
2 0 7 0 0 0 0 9 0 0 20 2
201 300
201 306
1 3 11 0 0 8320 0 7 9 0 0 3
101 219
101 222
169 222
1 0 3 0 0 0 0 6 0 0 21 2
135 69
135 128
1 0 4 0 0 0 0 8 0 0 22 2
92 72
92 107
0 0 2 0 0 4224 0 0 0 0 0 2
88 480
978 480
0 0 8 0 0 4224 0 0 0 0 0 2
82 335
981 335
0 0 7 0 0 4224 0 0 0 0 0 2
78 306
982 306
0 0 3 0 0 4224 0 0 0 0 0 2
67 128
982 128
0 0 4 0 0 4224 0 0 0 0 0 2
64 107
983 107
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
978 465 1007 489
988 473 996 489
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
982 321 1019 345
992 329 1008 345
2 M1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
985 290 1022 314
995 298 1011 314
2 M0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
983 111 1020 135
993 119 1009 135
2 I1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
984 90 1021 114
994 98 1010 114
2 I0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
