CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
-1424 28 -2 779
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
74 C:\Users\Lagoa\OneDrive\�rea de Trabalho\pes\projetos\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
-1256 124 -1143 221
9961490 0
0
6 Title:
5 Name:
0
0
0
26
12 IAGO.Mux.4x1
94 184 747 0 1 15
0 0
12 IAGO.Mux.4x1
17 0 4224 0
0
2 U8
71 3 85 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3820 0 0
2
45190.7 295
0
11 IAGO.Add.4b
94 860 244 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
11 IAGO.Add.4b
16 0 4224 0
0
2 U7
77 1 91 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7678 0 0
2
45190.7 225
0
13 IAGO.Buffer.4
94 676 245 0 8 17
0 14 15 17 16 10 11 12 13
13 IAGO.Buffer.4
15 0 4224 0
0
2 U6
76 0 90 8
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
961 0 0
2
45190.7 210
0
12 IAGO.Nand.4b
94 479 241 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
12 IAGO.Nand.4b
14 0 4224 0
0
2 U5
87 -2 101 6
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3178 0 0
2
45190.7 190
0
11 IAGO.Sub.4b
94 297 238 0 12 25
0 14 15 16 17 10 11 12 13 6
7 8 9
11 IAGO.Sub.4b
13 0 4224 0
0
2 U4
80 2 94 10
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3409 0 0
2
45190.7 120
0
14 Logic Display~
6 845 52 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
45190.7 119
0
14 Logic Display~
6 823 53 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
45190.7 118
0
14 Logic Display~
6 797 52 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
45190.7 117
0
14 Logic Display~
6 775 53 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
45190.7 116
0
8 Hex Key~
166 732 52 0 11 12
0 13 12 11 10 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9442 0 0
2
45190.7 115
0
8 Hex Key~
166 930 58 0 11 12
0 9 8 7 6 0 0 0 0 0
12 67
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9424 0 0
2
45190.7 114
0
14 Logic Display~
6 1058 48 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
45190.7 113
0
14 Logic Display~
6 1033 49 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
45190.7 112
0
14 Logic Display~
6 1009 49 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
45190.7 111
0
14 Logic Display~
6 987 49 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
45190.7 110
0
14 Logic Display~
6 1069 782 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
45190.7 109
0
14 Logic Display~
6 1094 782 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
45190.7 108
0
14 Logic Display~
6 1119 782 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
45190.7 107
0
14 Logic Display~
6 1141 781 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 U0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
45190.7 106
0
12 Hex Display~
7 1019 791 0 16 19
10 17 16 15 14 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
4 BusU
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6874 0 0
2
45190.7 105
0
12 IAGO.Mux.4x1
94 369 749 0 1 15
0 0
12 IAGO.Mux.4x1
12 0 4224 0
0
2 U9
71 3 85 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
5305 0 0
2
45190.7 71
0
12 IAGO.Mux.4x1
94 563 749 0 1 15
0 0
12 IAGO.Mux.4x1
11 0 4224 0
0
3 U10
68 3 89 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
34 0 0
2
45190.7 37
0
12 IAGO.Mux.4x1
94 744 750 0 1 15
0 0
12 IAGO.Mux.4x1
10 0 4224 0
0
3 U11
68 3 89 11
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
969 0 0
2
45190.7 3
0
8 Hex Key~
166 926 745 0 11 12
0 13 12 11 10 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 Ctrl
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8402 0 0
2
45190.7 2
0
14 Logic Display~
6 953 753 0 1 2
10 0
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
45190.7 1
0
14 Logic Display~
6 974 752 0 1 2
10 0
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
45190.7 0
0
135
2 0 0 0 0 272 0 23 0 0 15 3
666 772
655 772
655 823
1 0 0 0 0 272 0 23 0 0 16 3
666 750
651 750
651 812
2 0 0 0 0 272 0 22 0 0 15 3
485 771
473 771
473 823
1 0 0 0 0 272 0 22 0 0 16 3
485 749
466 749
466 812
2 0 0 0 0 272 0 21 0 0 15 3
291 771
284 771
284 823
1 0 0 0 0 272 0 21 0 0 16 3
291 749
278 749
278 812
7 0 0 0 0 16 0 23 0 0 65 2
744 794
744 837
7 0 0 0 0 16 0 22 0 0 64 2
563 793
563 845
7 0 0 0 0 16 0 21 0 0 63 2
369 793
369 856
7 0 0 0 0 16 0 1 0 0 62 2
184 791
184 864
2 0 0 0 0 16 0 24 0 0 15 2
929 769
929 823
1 0 0 0 0 16 0 24 0 0 16 2
935 769
935 812
1 0 0 0 0 272 0 25 0 0 15 2
953 771
953 823
1 0 0 0 0 272 0 26 0 0 16 2
974 770
974 812
2 0 0 0 0 272 0 1 0 0 0 4
106 769
101 769
101 823
987 823
1 0 0 0 0 272 0 1 0 0 0 4
106 747
98 747
98 812
987 812
6 0 0 0 0 16 0 22 0 0 76 2
570 719
570 498
3 0 0 0 0 16 0 23 0 0 69 2
693 719
693 635
4 0 0 0 0 16 0 23 0 0 73 2
724 721
724 560
6 0 0 0 0 16 0 23 0 0 77 2
751 720
751 481
5 0 0 0 0 16 0 23 0 0 81 2
777 720
777 411
4 0 0 0 0 16 0 22 0 0 71 2
543 720
543 589
3 0 0 0 0 16 0 22 0 0 68 2
512 718
512 652
5 0 0 0 0 16 0 22 0 0 80 2
596 719
596 428
3 0 0 0 0 16 0 21 0 0 67 2
318 718
318 664
4 0 0 0 0 16 0 21 0 0 72 2
349 720
349 577
6 0 0 0 0 16 0 21 0 0 76 2
376 719
376 498
5 0 0 0 0 16 0 21 0 0 79 2
402 719
402 440
3 0 0 0 0 16 0 1 0 0 66 2
133 716
133 677
4 0 0 0 0 16 0 1 0 0 70 2
164 718
164 602
6 0 0 0 0 16 0 1 0 0 74 2
191 717
191 523
5 0 0 0 0 16 0 1 0 0 78 2
217 717
217 453
1 0 0 0 0 16 0 5 0 0 66 2
261 284
261 677
2 0 0 0 0 16 0 5 0 0 67 2
288 282
288 664
3 0 0 0 0 16 0 5 0 0 68 2
315 284
315 652
4 0 0 0 0 16 0 5 0 0 69 2
343 283
343 635
1 0 0 0 0 16 0 4 0 0 70 2
439 288
439 602
2 0 0 0 0 16 0 4 0 0 71 2
467 288
467 589
3 0 0 0 0 16 0 4 0 0 72 2
502 289
502 577
4 0 0 0 0 16 0 4 0 0 73 2
538 288
538 560
1 0 0 0 0 16 0 3 0 0 74 2
631 284
631 523
2 0 0 0 0 16 0 3 0 0 75 2
656 285
656 510
4 0 0 0 0 16 0 3 0 0 76 2
685 284
685 498
3 0 0 0 0 16 0 3 0 0 77 2
713 283
713 481
1 0 0 0 0 16 0 2 0 0 78 2
824 289
824 453
2 0 0 0 0 16 0 2 0 0 79 2
851 289
851 440
3 0 0 0 0 16 0 2 0 0 80 2
878 288
878 428
4 0 0 0 0 16 0 2 0 0 81 2
905 288
905 411
0 0 0 0 0 272 0 0 0 0 0 5
1090 625
1090 688
1158 688
1158 625
1090 625
0 0 0 0 0 272 0 0 0 0 0 5
1090 553
1090 614
1157 614
1157 553
1090 553
0 0 0 0 0 272 0 0 0 0 0 5
1088 537
1088 475
1157 475
1157 541
1088 541
0 0 0 0 0 272 0 0 0 0 0 5
1084 374
1084 466
1155 466
1155 374
1084 374
0 0 3 0 0 272 0 0 0 0 0 8
1151 878
1151 829
1195 829
1195 889
1149 889
1149 875
1151 875
1151 874
4 0 14 0 0 16 0 20 0 0 62 2
1010 815
1010 864
3 0 15 0 0 16 0 20 0 0 63 2
1016 815
1016 856
2 0 16 0 0 16 0 20 0 0 64 2
1022 815
1022 845
1 0 17 0 0 16 0 20 0 0 65 2
1028 815
1028 837
1 0 14 0 0 16 0 16 0 0 62 2
1069 800
1069 864
1 0 15 0 0 16 0 17 0 0 63 2
1094 800
1094 856
1 0 16 0 0 16 0 18 0 0 64 2
1119 800
1119 845
1 0 17 0 0 16 0 19 0 0 65 2
1141 799
1141 837
0 0 14 0 0 16 0 0 0 0 0 2
99 864
1155 864
0 0 15 0 0 16 0 0 0 0 0 2
98 856
1156 856
0 0 16 0 0 16 0 0 0 0 0 2
98 845
1154 845
0 0 17 0 0 16 0 0 0 0 0 2
97 837
1155 837
0 0 0 0 0 16 0 0 0 0 0 2
93 677
1135 677
0 0 0 0 0 16 0 0 0 0 0 2
90 664
1136 664
0 0 0 0 0 16 0 0 0 0 0 2
89 652
1136 652
0 0 0 0 0 16 0 0 0 0 0 2
89 635
1137 635
0 0 0 0 0 16 0 0 0 0 0 2
91 602
1133 602
0 0 0 0 0 16 0 0 0 0 0 2
88 589
1134 589
0 0 0 0 0 16 0 0 0 0 0 2
87 577
1134 577
0 0 0 0 0 16 0 0 0 0 0 2
87 560
1135 560
0 0 0 0 0 16 0 0 0 0 0 2
90 523
1132 523
0 0 0 0 0 16 0 0 0 0 0 2
87 510
1133 510
0 0 0 0 0 16 0 0 0 0 0 2
86 498
1133 498
0 0 0 0 0 16 0 0 0 0 0 2
86 481
1134 481
0 0 0 0 0 16 0 0 0 0 0 2
91 453
1133 453
0 0 0 0 0 16 0 0 0 0 0 2
88 440
1134 440
0 0 0 0 0 16 0 0 0 0 0 2
87 428
1134 428
0 0 0 0 0 16 0 0 0 0 0 2
87 411
1135 411
0 0 4 0 0 272 0 0 0 0 0 5
1131 179
1131 137
1162 137
1162 179
1131 179
0 0 5 0 0 272 0 0 0 0 0 7
1121 71
1121 126
1155 126
1155 68
1122 68
1122 71
1121 71
9 0 6 0 0 16 0 2 0 0 120 2
883 211
883 171
10 0 7 0 0 16 0 2 0 0 121 2
893 210
893 163
11 0 8 0 0 16 0 2 0 0 122 2
901 210
901 152
12 0 9 0 0 16 0 2 0 0 123 2
911 211
911 144
5 0 10 0 0 16 0 2 0 0 132 2
810 211
810 116
6 0 11 0 0 16 0 2 0 0 133 2
820 211
820 108
7 0 12 0 0 16 0 2 0 0 134 2
830 211
830 97
8 0 13 0 0 16 0 2 0 0 135 2
839 211
839 89
5 0 10 0 0 16 0 3 0 0 132 2
631 210
631 116
6 0 11 0 0 16 0 3 0 0 133 2
658 210
658 108
7 0 12 0 0 16 0 3 0 0 134 2
685 212
685 97
8 0 13 0 0 16 0 3 0 0 135 2
714 211
714 89
9 0 6 0 0 16 0 4 0 0 120 2
507 198
507 171
10 0 7 0 0 16 0 4 0 0 121 2
520 198
520 163
11 0 8 0 0 16 0 4 0 0 122 2
535 198
535 152
12 0 9 0 0 16 0 4 0 0 123 2
546 199
546 144
5 0 10 0 0 16 0 4 0 0 132 2
426 199
426 116
6 0 11 0 0 16 0 4 0 0 133 2
444 198
444 108
7 0 12 0 0 16 0 4 0 0 134 2
462 198
462 97
8 0 13 0 0 16 0 4 0 0 135 2
479 198
479 89
9 0 6 0 0 16 0 5 0 0 120 2
324 204
324 171
10 0 7 0 0 16 0 5 0 0 121 2
333 204
333 163
11 0 8 0 0 16 0 5 0 0 122 2
342 203
342 152
12 0 9 0 0 16 0 5 0 0 123 2
352 204
352 144
5 0 10 0 0 16 0 5 0 0 132 2
244 204
244 116
6 0 11 0 0 16 0 5 0 0 133 2
257 205
257 108
7 0 12 0 0 16 0 5 0 0 134 2
270 204
270 97
8 0 13 0 0 16 0 5 0 0 135 2
279 204
279 89
4 0 6 0 0 16 0 11 0 0 120 2
921 82
921 171
3 0 7 0 0 16 0 11 0 0 121 2
927 82
927 163
2 0 8 0 0 16 0 11 0 0 122 2
933 82
933 152
1 0 9 0 0 16 0 11 0 0 123 2
939 82
939 144
1 0 6 0 0 16 0 15 0 0 120 2
987 67
987 171
1 0 7 0 0 16 0 14 0 0 121 2
1009 67
1009 163
1 0 8 0 0 16 0 13 0 0 122 2
1033 67
1033 152
1 0 9 0 0 16 0 12 0 0 123 2
1058 66
1058 144
0 0 6 0 0 16 0 0 0 0 0 2
84 171
1140 171
0 0 7 0 0 16 0 0 0 0 0 2
83 163
1141 163
0 0 8 0 0 16 0 0 0 0 0 2
83 152
1139 152
0 0 9 0 0 16 0 0 0 0 0 2
82 144
1140 144
4 0 10 0 0 16 0 10 0 0 132 2
723 76
723 116
3 0 11 0 0 16 0 10 0 0 133 2
729 76
729 108
2 0 12 0 0 16 0 10 0 0 134 2
735 76
735 97
1 0 13 0 0 16 0 10 0 0 135 2
741 76
741 89
1 0 10 0 0 16 0 9 0 0 132 2
775 71
775 116
1 0 11 0 0 16 0 8 0 0 133 2
797 70
797 108
1 0 12 0 0 16 0 7 0 0 134 2
823 71
823 97
1 0 13 0 0 16 0 6 0 0 135 2
845 70
845 89
0 0 10 0 0 16 0 0 0 0 0 2
80 116
1136 116
0 0 11 0 0 16 0 0 0 0 0 2
79 108
1137 108
0 0 12 0 0 16 0 0 0 0 0 2
79 97
1135 97
0 0 13 0 0 16 0 0 0 0 0 2
78 89
1136 89
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
853 15 906 39
863 23 895 39
4 IN'S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1162 143 1215 167
1172 151 1204 167
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1158 79 1211 103
1168 87 1200 103
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1193 843 1246 867
1203 851 1235 867
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1071 725 1116 749
1081 733 1105 749
3 OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1174 637 1227 661
1184 645 1216 661
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1179 654 1224 678
1189 662 1213 678
3 Sub
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1170 553 1223 577
1180 561 1212 577
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1171 569 1224 593
1181 577 1213 593
4 Nand
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1169 474 1222 498
1179 482 1211 498
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1163 491 1232 515
1173 499 1221 515
6 Buffer
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1171 400 1224 424
1181 408 1213 424
4 BusW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1173 418 1218 442
1183 426 1207 442
3 Add
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
905 683 982 707
915 691 971 707
7 Fun��es
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
