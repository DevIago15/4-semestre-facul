CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
61 C:\Users\Lagoa\OneDrive\�rea de Trabalho\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
14 Logic Display~
6 334 157 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5130 0 0
2
45185.7 0
0
14 Logic Display~
6 354 157 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
45185.7 1
0
14 Logic Display~
6 374 158 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
45185.7 2
0
9 2-In XOR~
219 406 278 0 3 22
0 6 5 9
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 XO1B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3421 0 0
2
45185.7 3
0
14 Logic Display~
6 644 158 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
45185.7 4
0
14 Logic Display~
6 665 157 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 W
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
45185.7 5
0
9 2-In XOR~
219 497 235 0 3 22
0 4 9 3
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 XO1A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
45185.7 6
0
9 2-In AND~
219 411 359 0 3 22
0 6 5 7
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 AN1B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7361 0 0
2
45185.7 7
0
9 2-In AND~
219 498 316 0 3 22
0 9 4 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 AN1A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
45185.7 8
0
8 2-In OR~
219 583 355 0 3 22
0 8 7 2
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 O1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
45185.7 9
0
8 Hex Key~
166 277 177 0 11 12
0 4 5 6 13 0 0 0 0 0
3 51
0
0 0 4656 0
0
6 SOURCE
-21 -34 21 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3472 0 0
2
45185.7 10
0
12 Hex Display~
7 727 186 0 18 19
10 3 2 14 15 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
7 DECIMAL
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9998 0 0
2
45185.7 11
0
11 IAGO.Add.1b
94 497 490 0 5 11
0 3 6 5 2 4
11 IAGO.Add.1b
1 0 4240 0
0
2 U1
70 -40 84 -32
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.90093e-315 0
0
34
4 0 2 0 0 8320 0 13 0 0 6 3
420 490
420 555
644 555
1 0 3 0 0 8192 0 13 0 0 7 3
497 524
497 532
665 532
0 5 4 0 0 4096 0 0 13 8 0 3
374 424
565 424
565 494
0 3 5 0 0 4096 0 0 13 9 0 3
354 429
542 429
542 457
0 2 6 0 0 4096 0 0 13 10 0 3
334 433
442 433
442 457
0 0 2 0 0 0 0 0 0 31 0 2
644 395
644 573
0 0 3 0 0 4096 0 0 0 30 0 2
665 395
665 574
0 0 4 0 0 0 0 0 0 32 0 2
374 393
374 574
0 0 5 0 0 0 0 0 0 33 0 2
354 394
354 575
0 0 6 0 0 4096 0 0 0 34 0 2
334 391
334 575
2 0 2 0 0 0 0 12 0 0 31 3
730 210
730 223
644 223
1 0 3 0 0 0 0 12 0 0 30 3
736 210
736 215
665 215
3 0 6 0 0 0 0 11 0 0 34 3
274 201
274 223
334 223
2 0 5 0 0 0 0 11 0 0 33 3
280 201
280 213
354 213
1 0 4 0 0 0 0 11 0 0 32 2
286 201
374 201
0 0 6 0 0 4480 0 0 0 0 0 6
318 179
678 179
678 399
320 399
320 179
322 179
3 2 7 0 0 4224 0 8 10 0 0 4
432 359
534 359
534 364
570 364
3 0 2 0 0 0 0 10 0 0 31 2
616 355
644 355
3 1 8 0 0 4224 0 9 10 0 0 4
519 316
550 316
550 346
570 346
2 0 4 0 0 0 0 9 0 0 32 2
474 325
374 325
1 0 9 0 0 4096 0 9 0 0 22 2
474 307
452 307
0 0 9 0 0 4352 0 0 0 27 0 2
452 278
452 311
2 0 5 0 0 0 0 8 0 0 33 2
387 368
354 368
1 0 6 0 0 0 0 8 0 0 34 2
387 350
334 350
3 0 3 0 0 0 0 7 0 0 30 2
530 235
665 235
1 0 4 0 0 0 0 7 0 0 32 2
481 226
374 226
3 2 9 0 0 8320 0 4 7 0 0 4
439 278
454 278
454 244
481 244
2 0 5 0 0 0 0 4 0 0 33 2
390 287
354 287
1 0 6 0 0 0 0 4 0 0 34 2
390 269
334 269
1 0 3 0 0 4224 0 6 0 0 0 2
665 175
665 400
1 0 2 0 0 0 0 5 0 0 0 2
644 176
644 400
1 0 4 0 0 4224 0 3 0 0 0 2
374 176
374 400
1 0 5 0 0 4224 0 2 0 0 0 2
354 175
354 400
1 0 6 0 0 0 0 1 0 0 16 2
334 175
334 399
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
447 137 540 161
457 145 529 161
9 Add. 1bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
572 177 609 201
582 185 598 201
2 L3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
500 176 537 200
510 184 526 200
2 L2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
403 174 440 198
413 182 429 198
2 L1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
